// Verilog netlist created by Tang Dynasty v5.5.47752
// Wed Jun 15 20:35:30 2022

`timescale 1ns / 1ps
module TEMAC_CORE
  (
  gmii_col,
  gmii_crs,
  gmii_rx_er,
  gmii_rx_vld,
  gmii_rxd,
  gmii_tx_clken,
  mac_cfg_vector,
  mdio_in,
  pause_req,
  pause_source_addr,
  pause_val,
  reset,
  rx_clk_en,
  rx_mac_clk,
  s_axi_aclk,
  s_axi_araddr,
  s_axi_arvalid,
  s_axi_awaddr,
  s_axi_awvalid,
  s_axi_bready,
  s_axi_rready,
  s_axi_wdata,
  s_axi_wvalid,
  tx_clk_en,
  tx_data,
  tx_data_en,
  tx_ifg_val,
  tx_mac_clk,
  tx_stop,
  unicast_addr,
  gmii_tx_en,
  gmii_tx_er,
  gmii_txd,
  mdio_clk,
  mdio_oen,
  mdio_out,
  rx_correct_frame,
  rx_data,
  rx_data_vld,
  rx_error_frame,
  rx_status_vector,
  rx_status_vld,
  s_axi_arready,
  s_axi_awready,
  s_axi_bresp,
  s_axi_bvalid,
  s_axi_rdata,
  s_axi_rresp,
  s_axi_rvalid,
  s_axi_wready,
  speed_10,
  speed_100,
  speed_1000,
  tx_collision,
  tx_rdy,
  tx_retransmit,
  tx_status_vector,
  tx_status_vld
  );

  input gmii_col;
  input gmii_crs;
  input gmii_rx_er;
  input gmii_rx_vld;
  input [7:0] gmii_rxd;
  input gmii_tx_clken;
  input [19:0] mac_cfg_vector;
  input mdio_in;
  input pause_req;
  input [47:0] pause_source_addr;
  input [15:0] pause_val;
  input reset;
  input rx_clk_en;
  input rx_mac_clk;
  input s_axi_aclk;
  input [7:0] s_axi_araddr;
  input s_axi_arvalid;
  input [7:0] s_axi_awaddr;
  input s_axi_awvalid;
  input s_axi_bready;
  input s_axi_rready;
  input [31:0] s_axi_wdata;
  input s_axi_wvalid;
  input tx_clk_en;
  input [7:0] tx_data;
  input tx_data_en;
  input [7:0] tx_ifg_val;
  input tx_mac_clk;
  input tx_stop;
  input [47:0] unicast_addr;
  output gmii_tx_en;
  output gmii_tx_er;
  output [7:0] gmii_txd;
  output mdio_clk;
  output mdio_oen;
  output mdio_out;
  output rx_correct_frame;
  output [7:0] rx_data;
  output rx_data_vld;
  output rx_error_frame;
  output [26:0] rx_status_vector;
  output rx_status_vld;
  output s_axi_arready;
  output s_axi_awready;
  output [1:0] s_axi_bresp;
  output s_axi_bvalid;
  output [31:0] s_axi_rdata;
  output [1:0] s_axi_rresp;
  output s_axi_rvalid;
  output s_axi_wready;
  output speed_10;
  output speed_100;
  output speed_1000;
  output tx_collision;
  output tx_rdy;
  output tx_retransmit;
  output [28:0] tx_status_vector;
  output tx_status_vld;

  parameter P_ADD_FILT_EN = 1'b1;
  parameter P_ADD_FILT_LIST = 3;
  parameter P_HALF_DUPLEX = 1'b1;
  parameter P_HOST_EN = 1'b1;
  parameter P_SPEED_1000 = 1'b0;
  parameter P_SPEED_10_100 = 1'b0;
  parameter P_TRI_SPEED = 1'b1;
  // localparam P_CLK_EN = 1'b1;
  wire [15:0] al_2c28b3bd;
  wire [15:0] al_a6672453;
  wire [4:0] al_bd4c52f0;
  wire [7:0] al_e8c856c9;
  wire [4:0] al_d002eac;
  wire [15:0] al_b9f27169;
  wire [7:0] al_45ed4524;
  wire [4:0] al_1dee2dce;
  wire [47:0] al_9fdb6cdc;
  wire [15:0] al_27d2fc1a;
  wire [2:0] al_d97145b1;
  wire  al_14405a50;
  wire  al_36ab2fb9;
  wire  al_e61a7e67;
  wire  al_b47e09b3;
  wire  al_91e39671;
  wire  al_88c8ee13;
  wire  al_b8dbdfec;
  wire  al_7bcff3b9;
  wire  al_9d9cd237;
  wire  al_ed22e70c;
  wire  al_83ef8a4e;
  wire [4:0] al_7c53cb60;
  wire [7:0] al_9c572362;
  wire [7:0] al_251fb86c;
  wire [15:0] al_ac3dcbf8;
  wire [5:0] al_38c57749;
  wire [5:0] al_9868190b;
  wire [15:0] al_dd86ad38;
  wire [15:0] al_a128253b;
  wire [14:0] al_b79f6a7b;
  wire [7:0] al_ecbdcaf1;
  wire [3:0] al_2e624116;
  wire [3:0] al_d286f1cd;
  wire [3:0] al_62f364a9;
  wire [7:0] al_fbc4ef28;
  wire [11:0] al_d2863baf;
  wire [3:0] al_a59c7c46;
  wire [3:0] al_20d4193c;
  wire [3:0] al_96252128;
  wire [7:0] al_b25edb3;
  wire [7:0] al_78b1b46e;
  wire [7:0] al_5bef7ee6;
  wire [3:0] al_dc435ff2;
  wire [3:0] al_ee96b553;
  wire [3:0] al_95650af7;
  wire [7:0] al_fa90a029;
  wire [7:0] al_bb772f98;
  wire [7:0] al_5160c8c2;
  wire [7:0] al_5db4ba74;
  wire [5:0] al_ddeffb0f;
  wire [5:0] al_58820abe;
  wire [15:0] al_89a4ecab;
  wire [7:0] al_82716c38;
  wire [7:0] al_13660933;
  wire [31:0] al_88fb5330;
  wire [31:0] al_7808e039;
  wire [6:0] al_4096d0c7;
  wire [31:0] al_523025ae;
  wire [31:0] al_ab2a7f1;
  wire [31:0] al_238a702c;
  wire [31:0] al_939ca227;
  wire [7:0] al_3833d624;
  wire [7:0] al_7b2ceef0;
  wire [31:0] al_492d1bb8;
  wire [31:0] al_868a1cad;
  wire [31:0] al_cd0aa0ee;
  wire [31:0] al_a0f12bef;
  wire  al_f3899d20;
  wire [1:0] al_25215c55;
  wire [31:0] al_9b4eaefc;
  wire  al_4db525a4;
  wire  al_c3f8fcfd;
  wire  al_62e089bb;
  wire  al_33409841;
  wire  al_eb828cf9;
  wire  al_53937ca8;
  wire  al_75328a30;
  wire  al_6bda5d58;
  wire  al_47962165;
  wire [5:0] al_ec1f16c4;
  wire [15:0] al_9f0e53e2;
  wire [15:0] al_8867ef3c;
  wire [15:0] al_628888c;
  wire [31:0] al_39eeae1d;
  wire [3:0] al_5ea2be94;
  wire [31:0] al_220ff640;
  wire [9:0] al_be957c85;
  wire [9:0] al_aea26701;
  wire [9:0] al_1ac19429;
  wire [15:0] al_aac09418;
  wire [14:0] al_cbc62139;
  wire [15:0] al_14016c23;
  wire [1:0] al_d6a2be89;
  wire [14:0] al_c86ca47d;
  wire [14:0] al_92477e6d;
  wire [15:0] al_f0afd253;
  wire [15:0] al_73eb08b7;
  wire [7:0] al_e8c5f626;
  wire [7:0] al_4b3fffb5;
  wire [7:0] al_b242ee60;
  wire [7:0] al_12d2a17a;
  wire [5:0] al_54f03dbf;
  wire [1:0] al_71b48cc2;
  wire [3:0] al_516522f9;
  wire [13:0] al_1f0d50be;
  wire [24:0] al_c5802d0a;
  wire [1:0] al_b1b61f7c;
  wire [15:0] al_ba4af77d;
  wire [15:0] al_93bf05b4;
  wire [15:0] al_4c524efc;
  wire [15:0] al_f4c47e2b;
  wire [15:0] al_5d5249da;
  wire [15:0] al_f6dc28d8;
  wire [15:0] al_d5e21796;
  wire [15:0] al_d57700f8;
  wire [9:0] al_6c9db937;
  wire [14:0] al_ae5f998b;
  wire [13:0] al_e1759dc;
  wire [3:0] al_ed1f021e;
  wire [2:0] al_e702d1c;
  wire [3:0] al_3a9d8027;
  wire [2:0] al_536d34;
  wire [12:0] al_715819dc;
  wire [1:0] al_b01f953d;
  wire [13:0] al_72a2cf60;
  wire [1:0] al_ed15c12c;
  wire [12:0] al_1f1bbfc9;
  wire [9:0] al_6e9a1ae;
  wire [3:0] al_e23c1f65;
  wire [5:0] al_5f257019;
  wire [18:0] al_e8bb9040;
  wire [14:0] al_efc7f78a;
  wire [14:0] al_64fd2ef5;
  wire [14:0] al_183e87f4;
  wire [31:0] al_2cf31306;
  wire [3:0] al_b130642e;
  wire [31:0] al_a7d56e64;
  wire [1:0] al_77f0ddfc;
  wire [7:0] al_4d46dbf7;
  wire [7:0] al_9affd881;
  wire [7:0] al_84c0beb4;
  wire [7:0] al_8a6ca59e;
  wire [7:0] al_e00c8785;
  wire [7:0] al_96e5a141;
  wire [14:0] al_8e462c61;
  wire [10:0] al_8c490204;
  wire [14:0] al_e512aff;
  wire [14:0] al_19bf88c2;
  wire [7:0] al_54d2aa3;
  wire [13:0] al_24da7d44;
  wire [7:0] al_984d3b84;
  wire [7:0] al_67d6ec64;
  wire [3:0] al_bef8ea23;
  wire [1:0] al_f3f63e4d;
  wire [9:0] al_821706b3;
  wire [15:0] al_bff87853;
  wire [13:0] al_48fcd383;
  wire [2:0] al_24ac8493;
  wire [1:0] al_e4dc5a7;
  wire [7:0] al_84a48183;
  wire [2:0] al_63a836a9;
  wire [7:0] al_6ec37834;
  wire [7:0] al_c122424e;
  wire [1:0] al_b3968bab;
  wire [1:0] al_630a3426;
  wire [19:0] al_acbf9207;
  wire [18:0] al_77695f5b;
  wire [5:0] al_20b55994;
  wire [14:0] al_f5f472e;
  wire [14:0] al_c007c6a1;
  wire [4:0] al_ae339d26;
  wire [7:0] al_224d6023;
  wire [7:0] al_93cc3d71;
  wire [7:0] al_9595c97a;
  wire [7:0] al_f83013e9;
  wire [14:0] al_ecab3deb;
  wire [15:0] al_e20fd0c7;
  wire [14:0] al_4b4b7bbc;
  wire [9:0] al_dcce7f97;
  wire [9:0] al_93f1315e;
  wire [10:0] al_c8474427;
  wire [63:0] al_752f7592;
  wire [63:0] al_d1b76c6b;
  wire [63:0] al_902efd00;
  wire [3:0] al_b9297703;
  wire [2:0] al_d0555e9d;
  wire [15:0] al_ecfcb422;
  wire [127:0] al_3a736cff;
  wire  al_e7f17f52;
  wire  al_e774f130;
  wire  al_7ce61a6c;
  wire  al_b292fc1;
  wire  al_9e1e2a36;
  wire  al_8fcbb835;
  wire  al_6e6c13e6;
  wire  al_c9f27122;
  wire  al_3a099803;
  wire  al_1d49aa78;
  wire  al_67882c63;
  wire  al_133f55a2;
  wire  al_d849110a;
  wire  al_f8a9808f;
  wire  al_50c6f567;
  wire  al_95dcd5c9;
  wire  al_d9e64745;
  wire  al_47ed325a;
  wire  al_67edee18;
  wire  al_3255583f;
  wire  al_b91e0498;
  wire  al_ec16c3b2;
  wire  al_71c12aaa;
  wire  al_2f3d50c1;
  wire  al_65907c46;
  wire  al_5c5a5e75;
  wire  al_c7b03fcb;
  wire  al_70936044;
  wire  al_5e3e1251;
  wire  al_a51c3dde;
  wire  al_29fafdbd;
  wire  al_2cc28140;
  wire [31:0] al_e6b493f;
  wire [47:0] al_40f6174;
  wire [47:0] al_f0cac652;
  wire [47:0] al_9db0b0fa;
  wire [2:0] al_7e8a07be;
  wire [47:0] al_2408f449;
  wire  al_a4fb2b45;
  wire  al_6a6bba48;
  wire  al_c3e9514;
  wire  al_f1396ae3;
  wire  al_da9f8ded;
  wire  al_655153ec;
  wire  al_8ba02654;
  wire  al_9993ad5e;
  wire  al_29e11b90;
  wire  al_d1a1cb58;
  wire  al_989215e7;
  wire  al_ac9336a;
  wire  al_9c616a92;
  wire  al_e19dcc16;
  wire  al_a4c57dd8;
  wire  al_e4b485d4;
  wire  al_a880ef2c;
  wire  al_1974d963;
  wire  al_b3009928;
  wire  al_f13bd74f;
  wire  al_2ad06c7e;
  wire  al_159c9d41;
  wire  al_fefd5fd3;
  wire  al_ca969cfa;
  wire  al_dd993167;
  wire  al_4285f2d3;
  wire  al_8b78b709;
  wire  al_c40403fa;
  wire  al_b6be24f;
  wire  al_ad7719c4;
  wire  al_eaf2c767;
  wire  al_8b492536;
  wire [7:0] al_5fe249d5;
  wire [47:0] al_49a90ce2;
  wire [47:0] al_2bdcc449;
  wire al_c58b187c;
  wire al_e6bb9c83;
  wire al_4c4d90b0;
  wire al_627de329;
  wire al_fc03cb77;
  wire al_63c928c0;
  wire al_c2c7d796;
  wire al_90021ccb;
  wire al_9f678f08;
  wire al_f6518188;
  wire al_737a8715;
  wire al_8765eb4;
  wire al_3fe33606;
  wire al_67074a64;
  wire al_87a09a9e;
  wire al_f03a2c10;
  wire al_1824196b;
  wire al_8b041f7e;
  wire al_e5699de4;
  wire al_70372a24;
  wire al_c00b2fb7;
  wire al_350ee797;
  wire al_e5314cad;
  wire al_64d29977;
  wire al_609ad6f2;
  wire al_70727c2f;
  wire al_8f322b4;
  wire al_11c159a;
  wire al_7cd2fee3;
  wire al_127a14bf;
  wire al_4dd161f2;
  wire al_179835d0;
  wire al_41b2f611;
  wire al_d7707346;
  wire al_3b505c23;
  wire al_ac5af120;
  wire al_d9170e3;
  wire al_61fb0a6;
  wire al_be16aa76;
  wire al_b2b8b63f;
  wire al_f4252f15;
  wire al_3aae9c28;
  wire al_346eaec2;
  wire al_644f021d;
  wire al_42966d4a;
  wire al_8c6ac38c;
  wire al_81681eb;
  wire al_18c1e35a;
  wire al_662270e8;
  wire al_a03de72f;
  wire al_9fbaf8f2;
  wire al_dbb71724;
  wire al_5006fa3b;
  wire al_53f52d8d;
  wire al_9fcf7528;
  wire al_4beb6793;
  wire al_acabe8fb;
  wire al_46ece34d;
  wire al_1caff122;
  wire al_826fce19;
  wire al_1d01387;
  wire al_8e145c1c;
  wire al_2c95779d;
  wire al_edb0b8cc;
  wire al_da9cd0a9;
  wire al_d8bac65b;
  wire al_438ac6ff;
  wire al_ca04b07a;
  wire al_2e8c1b28;
  wire al_68258153;
  wire al_a7af4189;
  wire al_32667361;
  wire al_ae33357f;
  wire al_67b92cd9;
  wire al_a9aea0ae;
  wire al_7a5b596f;
  wire al_ff9e33ad;
  wire al_591adfcf;
  wire al_5fd6768b;
  wire al_38ea72f1;
  wire al_810ba8de;
  wire al_8b51ab4;
  wire al_6ea32e9c;
  wire al_8b7d9749;
  wire al_8b780845;
  wire al_2337d80f;
  wire al_aa427d37;
  wire al_6d2cc211;
  wire al_1e2edecf;
  wire al_1a7bad30;
  wire al_e5091a32;
  wire al_46f5ce71;
  wire al_89fbca82;
  wire al_ed888342;
  wire al_88c53423;
  wire al_8399b753;
  wire al_7bec6b72;
  wire al_132ae268;
  wire al_e8564782;
  wire al_5df5c44f;
  wire al_72f5321b;
  wire al_61aea43e;
  wire al_9fe1548f;
  wire al_d3f3dfbd;
  wire al_2a91cf37;
  wire al_f13f5376;
  wire al_6b4499fc;
  wire al_fc3fb77f;
  wire al_e18a88b8;
  wire al_fcf500fb;
  wire al_7f87fb2e;
  wire al_ff9a7266;
  wire al_f517c689;
  wire al_59850dc4;
  wire al_90484227;
  wire al_f17b93eb;
  wire al_81344cef;
  wire al_6de80447;
  wire al_abc98a52;
  wire al_fc3c716f;
  wire al_7c94b9c5;
  wire al_e8fc825c;
  wire al_6b48ce98;
  wire al_77b8d1cd;
  wire al_59f1a9e9;
  wire al_ec74b2dd;
  wire al_dad1457e;
  wire al_2e1a2363;
  wire al_3fd53f68;
  wire al_1a6b1e5a;
  wire al_71becb96;
  wire al_2bb2d81d;
  wire al_678e4333;
  wire al_4f0de751;
  wire al_50f7b858;
  wire al_dc85d54;
  wire al_d61cd20b;
  wire al_7b7a3c37;
  wire al_5374577;
  wire al_ba2c5d76;
  wire al_a700dfa6;
  wire al_74b73e47;
  wire al_14acaf34;
  wire al_f7d4c035;
  wire al_92a04064;
  wire al_f6b6167;
  wire al_32868173;
  wire al_574485a3;
  wire al_8b27d348;
  wire al_98b546cc;
  wire al_2bf5454d;
  wire al_54e389b6;
  wire al_3956f95a;
  wire al_25ad8958;
  wire al_81b1fe1c;
  wire al_bde4ed05;
  wire al_6f2ddcc1;
  wire al_cde2200a;
  wire al_57e58431;
  wire al_776d5772;
  wire al_d293a382;
  wire al_be08372;
  wire al_4bb8f8b3;
  wire al_988cc37d;
  wire al_5f618b63;
  wire al_6219a09a;
  wire al_d4f64f24;
  wire al_bc58b1b4;
  wire al_bc147132;
  wire al_6e8a0941;
  wire al_b984f6c1;
  wire al_ee74aec5;
  wire al_77ced363;
  wire al_20c861d8;
  wire al_269c8a2f;
  wire al_c078e47f;
  wire al_c3d753a2;
  wire al_dbdc14b4;
  wire al_80471da6;
  wire al_f4dbb19c;
  wire al_6702ffbf;
  wire al_21291e01;
  wire al_5f71b9c1;
  wire al_b2ee3fbb;
  wire al_d5df3ac1;
  wire al_53bc66bd;
  wire al_d30618ea;
  wire al_9c3c5741;
  wire al_1c02a3cb;
  wire al_ae0d49cd;
  wire al_9df86c79;
  wire al_4f080ff4;
  wire al_f12d2a54;
  wire al_951148c8;
  wire al_3e63fd9;
  wire al_19dda09f;
  wire al_46b6d0af;
  wire al_20d13f12;
  wire al_3290811f;
  wire al_e25e65e3;
  wire al_607f31be;
  wire al_b5a71093;
  wire al_336a5970;
  wire al_700f8a99;
  wire al_633f8ef2;
  wire al_bc3d033e;
  wire al_89a3ef5a;
  wire al_b1d5fd9b;
  wire al_adcb0cbd;
  wire al_62884f47;
  wire al_b746bad7;
  wire al_27893604;
  wire al_c2dc89e9;
  wire al_7541e92c;
  wire al_6df60a04;
  wire al_e98fadb;
  wire al_8027e03;
  wire al_4e0a4dc5;
  wire al_d890a7e6;
  wire al_1ca8afe3;
  wire al_de12b3ef;
  wire al_dd6bc6a;
  wire al_87773c5e;
  wire al_c88c8301;
  wire al_29842798;
  wire al_68462158;
  wire al_3cd9a398;
  wire al_a09e8e00;
  wire al_cd1b7e74;
  wire al_b3be0d17;
  wire al_87969af9;
  wire al_7ac4c27f;
  wire al_8cc75feb;
  wire al_6b5283b3;
  wire al_10fc4c0e;
  wire al_54081406;
  wire al_dd9e938b;
  wire al_977227b4;
  wire al_fadd6423;
  wire al_520be21e;
  wire al_ec9f94d8;
  wire al_47e79db6;
  wire al_7868fcca;
  wire al_78567007;
  wire al_3efdaf7e;
  wire al_e4a226df;
  wire al_dbdccc1f;
  wire al_9bcb8f17;
  wire al_81191a79;
  wire al_a6edfc2;
  wire al_3abe5c64;
  wire al_f974815d;
  wire al_7f233c39;
  wire al_42136331;
  wire al_5832a18a;
  wire al_fde4e9e1;
  wire al_6b963607;
  wire al_e364ec9e;
  wire al_923f48aa;
  wire al_7b831e20;
  wire al_4d9c1d5;
  wire al_bc71f40f;
  wire al_1887f4c;
  wire al_ead880b8;
  wire al_57798083;
  wire al_64ec9565;
  wire al_4c385591;
  wire al_3fd7c40d;
  wire al_cf7c6c77;
  wire al_de861c69;
  wire al_bf96f833;
  wire al_191a34b5;
  wire al_8aa62a5b;
  wire al_3329776d;
  wire al_30bba5ae;
  wire al_f246f984;
  wire al_b8c67773;
  wire al_8319735a;
  wire al_639b4ff6;
  wire al_717e3e2b;
  wire al_8afbeabf;
  wire al_5c023966;
  wire al_44998c84;
  wire al_2179357c;
  wire al_5d1a6fb0;
  wire al_76966ac9;
  wire al_4f8a4577;
  wire al_ca9e38f4;
  wire al_f7494ece;
  wire al_bbe3a962;
  wire al_54fc2cdd;
  wire al_6300b493;
  wire al_65b028e9;
  wire al_c981d7f0;
  wire al_1ce38576;
  wire al_5f85f29c;
  wire al_d5243429;
  wire al_40a7c639;
  wire al_fbfd813b;
  wire al_ec490bfd;
  wire al_58bd59f6;
  wire al_ebd456eb;
  wire al_b59c2e50;
  wire al_575bbbae;
  wire al_6f9895cd;
  wire al_b0d2bfc8;
  wire al_73782b81;
  wire al_29cb65c6;
  wire al_7a2a1104;
  wire al_1e9fbff4;
  wire al_d2811bd8;
  wire al_f2cdbc14;
  wire al_fc353ce9;
  wire al_dfffc03a;
  wire al_f51408c3;
  wire al_5b8b9ce6;
  wire al_c91a5908;
  wire al_7fb47a00;
  wire al_1104f08c;
  wire al_ab14fdf9;
  wire al_25417591;
  wire al_ee8473c1;
  wire al_eeaafdd6;
  wire al_af3a6b91;
  wire al_d10bb6dd;
  wire al_95e117eb;
  wire al_361cbc23;
  wire al_dbee6318;
  wire al_36d5f4c5;
  wire al_fbb2ea7a;
  wire al_88a372db;
  wire al_a48c9e07;
  wire al_d0ab12fe;
  wire al_4f97dd8c;
  wire al_bb4cafc;
  wire al_9dbb5412;
  wire al_8e6b9688;
  wire al_aa5dc84f;
  wire al_96d069e8;
  wire al_68e39bd9;
  wire al_a140f198;
  wire al_900fca1b;
  wire al_d9ca5f64;
  wire al_cf085f09;
  wire al_3e886516;
  wire al_e199650d;
  wire al_6490a8fc;
  wire al_642e830e;
  wire al_643ac1f2;
  wire al_e3f5d0d6;
  wire al_f6643499;
  wire al_206f470e;
  wire al_8aa33695;
  wire al_1f250659;
  wire al_2a71f823;
  wire al_c925873;
  wire al_af6614da;
  wire al_ea441981;
  wire al_f731da11;
  wire al_d1e17be4;
  wire al_85bba154;
  wire al_fdd1f60e;
  wire al_c35ead5c;
  wire al_a494216e;
  wire al_1d8c2b07;
  wire al_4fb6999c;
  wire al_33f2071f;
  wire al_e1420a1f;
  wire al_f52ae365;
  wire al_177c7491;
  wire al_72403be8;
  wire al_6fa8f988;
  wire al_ee3bb963;
  wire al_548d2e8d;
  wire al_c52cf3e8;
  wire al_7fe117d0;
  wire al_12358921;
  wire al_5b769262;
  wire al_13f48428;
  wire al_56978088;
  wire al_6a534a0a;
  wire al_4d3e0511;
  wire al_c388f857;
  wire al_20a6f635;
  wire al_1f6fed00;
  wire al_bea385e7;
  wire al_d224660a;
  wire al_b7729dd8;
  wire al_7cd73f8f;
  wire al_eb5c4882;
  wire al_b348c1a2;
  wire al_e2a3cd9;
  wire al_e5fcf9b1;
  wire al_cbafc250;
  wire al_e396ca5d;
  wire al_d75651de;
  wire al_f2f960a1;
  wire al_2b1074ba;
  wire al_f92f3a06;
  wire al_d09ba8fa;
  wire al_21d722fe;
  wire al_b65fd623;
  wire al_567fa47e;
  wire al_f28e4921;
  wire al_64e175a6;
  wire al_4dac203f;
  wire al_8b86ece7;
  wire al_3475fb1c;
  wire al_6980bc30;
  wire al_1bfb1d64;
  wire al_af1ac2b6;
  wire al_75182ad3;
  wire al_5ad7d7e7;
  wire al_c5664b3b;
  wire al_9f6ea2ef;
  wire al_ad4aba0;
  wire al_d3482891;
  wire al_25d4a5f3;
  wire al_68ba43d4;
  wire al_9a8c459a;
  wire al_a978a29f;
  wire al_f92026f1;
  wire al_4b2213d6;
  wire al_edc29fee;
  wire al_d27166fa;
  wire al_c2463579;
  wire al_be1d3817;
  wire al_3620963e;
  wire al_b1328a1f;
  wire al_4a548f7c;
  wire al_ea30f787;
  wire al_77192586;
  wire al_1d84107f;
  wire al_5227328;
  wire al_1dbbddf2;
  wire al_af806095;
  wire al_97576f4d;
  wire al_64c768d;
  wire al_acdc1781;
  wire al_d6cf9565;
  wire al_ab89cd63;
  wire al_8640fd7b;
  wire al_df015ce6;
  wire al_f192c825;
  wire al_742c008b;
  wire al_29b24aa7;
  wire al_98e25f8d;
  wire al_9f207ad1;
  wire al_93b20b44;
  wire al_39bb46f4;
  wire al_a1a0ec14;
  wire al_f80c5908;
  wire al_17387d1;
  wire al_36605837;
  wire al_37f58acb;
  wire al_4421c6bd;
  wire al_acb6d76c;
  wire al_47b64b8f;
  wire al_4d7216c9;
  wire al_1698ebe9;
  wire al_3c6cc34f;
  wire al_1e340161;
  wire al_4be4ecdd;
  wire al_e04ba284;
  wire al_cf06a90;
  wire al_913e13a3;
  wire al_da8b063f;
  wire al_4f19e5d0;
  wire al_3b1a77d7;
  wire al_531ee03c;
  wire al_92cc5462;
  wire al_4973ef09;
  wire al_b62e571a;
  wire al_c59c6deb;
  wire al_638d20bb;
  wire al_8f030415;
  wire al_6b2f12fa;
  wire al_279c902b;
  wire al_51172105;
  wire al_8afe6a9f;
  wire al_952d11ed;
  wire al_24f8640d;
  wire al_69f453c2;
  wire al_a6c89001;
  wire al_81cdbd25;
  wire al_7ffb8465;
  wire al_ecd47e95;
  wire al_3557a617;
  wire al_e336c621;
  wire al_907f6029;
  wire al_2e2debcb;
  wire al_ccc3c4e3;
  wire al_34d2745e;
  wire al_b0eb70b2;
  wire al_5764731d;
  wire al_114ce5a4;
  wire al_4ba3ac36;
  wire al_a12adb97;
  wire al_4a89f542;
  wire al_70a59d2e;
  wire al_ffd3f5d1;
  wire al_a8d1cf64;
  wire al_1751a6d0;
  wire al_360cb20;
  wire al_eaacfd93;
  wire al_4fe9a477;
  wire al_bb3ef93c;
  wire al_8f22b7e0;
  wire al_cbbf04f9;
  wire al_1e8f68ca;
  wire al_75356484;
  wire al_1491ad5;
  wire al_db73eae9;
  wire al_aa6ddd9b;
  wire al_4e7d0870;
  wire al_964d579;
  wire al_397de144;
  wire al_32b11a18;
  wire al_b3c5207a;
  wire al_fa26b745;
  wire al_1a33f9b0;
  wire al_d277135;
  wire al_b156040b;
  wire al_f28fd6dc;
  wire al_7f7f4148;
  wire al_ab82ee9a;
  wire al_95d27a4c;
  wire al_8aeddbc;
  wire al_bca5d36c;
  wire al_7c03a443;
  wire al_8f0a5b42;
  wire al_cafc0d92;
  wire al_8b965f41;
  wire al_66382828;
  wire al_5156ba29;
  wire al_4854aa2f;
  wire al_e03ae0c1;
  wire al_5cd49131;
  wire al_508b6c4c;
  wire al_4d4a65fe;
  wire al_1638f286;
  wire al_44b2d585;
  wire al_6b4822fe;
  wire al_fc7de59c;
  wire al_f2d6f40b;
  wire al_3cdb7f2c;
  wire al_ee9e22e;
  wire al_addc1415;
  wire al_81aa4d04;
  wire al_756a1d77;
  wire al_54bdd1be;
  wire al_f4b18dcd;
  wire al_bfb14c0f;
  wire al_4c9c0764;
  wire al_275437c2;
  wire al_c78fe3c1;
  wire al_5411d218;
  wire al_e30f13e9;
  wire al_3d188dba;
  wire al_a7b91d29;
  wire al_219561f;
  wire al_4fb560ef;
  wire al_3d691a71;
  wire al_c9a41ba;
  wire al_eccfd98c;
  wire al_eefcdfd;
  wire al_58846bb5;
  wire al_6303158d;
  wire al_34d58259;
  wire al_69600a84;
  wire al_ebcb9742;
  wire al_7b06746d;
  wire al_bd268370;
  wire al_64206da8;
  wire al_922f69ff;
  wire al_baa25bac;
  wire al_22f4f2dd;
  wire al_7a3587c3;
  wire al_a162bb8e;
  wire al_3c42ccfe;
  wire al_46fe62ca;
  wire al_c504b787;
  wire al_beea368e;
  wire al_5ef35ad0;
  wire al_2c5269c;
  wire al_dc745a17;
  wire al_9b6b0ae2;
  wire al_f8bfe558;
  wire al_a49d6a86;
  wire al_4a547188;
  wire al_72ac780f;
  wire al_22c188eb;
  wire al_a6f148e9;
  wire al_674bc53d;
  wire al_26f70e9a;
  wire al_186c00a8;
  wire al_3c343df4;
  wire al_21c59f1;
  wire al_cd3fff34;
  wire al_52e770ef;
  wire al_5d53f279;
  wire al_7c904594;
  wire al_f785157a;
  wire al_3dc7e6d6;
  wire al_25dd3b31;
  wire al_8edce7a2;
  wire al_b4b52182;
  wire al_44e126e5;
  wire al_bb1dc6ea;
  wire al_7978050f;
  wire al_25291b5c;
  wire al_1cbba6e6;
  wire al_372f5c11;
  wire al_68634068;
  wire al_3119a20d;
  wire al_cb74bfe8;
  wire al_90c946f9;
  wire al_e202820f;
  wire al_c702b161;
  wire al_321e78bf;
  wire al_7bce675b;
  wire al_f9cac200;
  wire al_a7a7af9e;
  wire al_c2569e9f;
  wire al_d0a10128;
  wire al_3da78c22;
  wire al_db0897ce;
  wire al_603ec03;
  wire al_34784d5d;
  wire al_f16920e0;
  wire al_2f3f17d;
  wire al_6ecd5054;
  wire al_ce80051a;
  wire al_bbb4d320;
  wire al_391ec013;
  wire al_ed990b15;
  wire al_8e811a01;
  wire al_cd9c4b15;
  wire al_a14eea73;
  wire al_e4bdca8a;
  wire al_dc6fb7d9;
  wire al_32839ce1;
  wire al_316af0f0;
  wire al_ff67665e;
  wire al_531e5772;
  wire al_54d691ed;
  wire al_d632949b;
  wire al_cc4e6731;
  wire al_c5bc3747;
  wire al_d0ecc99e;
  wire al_49bc5cf4;
  wire al_9e8909aa;
  wire al_cac2565f;
  wire al_6c890ee8;
  wire al_d280e871;
  wire al_1feb4c09;
  wire al_e2b7a540;
  wire al_5772dfd3;
  wire al_43bf9cc4;
  wire al_921d9eff;
  wire al_da5fd7db;
  wire al_80344ab4;
  wire al_6baf9e53;
  wire al_749e1728;
  wire al_3252df70;
  wire al_7bee3de4;
  wire al_8d11b694;
  wire al_a87a1c23;
  wire al_6281ecee;
  wire al_f7f8cae;
  wire al_3e7ed8af;
  wire al_2ff03e70;
  wire al_d1ddae16;
  wire al_6627cbad;
  wire al_9907ae47;
  wire al_7701781b;
  wire al_d5b2f5c4;
  wire al_614db0a6;
  wire al_2e8ff7ab;
  wire al_77df94be;
  wire al_e06bfe23;
  wire al_535d21bf;
  wire al_b3eb9d64;
  wire al_289fe017;
  wire al_77be5888;
  wire al_7f375c7a;
  wire al_c1e4e3b;
  wire al_4b9a6e34;
  wire al_67caff7a;
  wire al_5ae0e8ee;
  wire al_6bfa7885;
  wire al_1a86743a;
  wire al_8f82c138;
  wire al_db547825;
  wire al_89eb3505;
  wire al_29f8870a;
  wire al_abc7ca1f;
  wire al_e8517c4;
  wire al_d1451a79;
  wire al_467061b3;
  wire al_b42812f4;
  wire al_38b760cc;
  wire al_7c0134d3;
  wire al_31ba2088;
  wire al_25b9a235;
  wire al_c9d3334;
  wire al_a021098c;
  wire al_e0f968c1;
  wire al_40bf3e87;
  wire al_baff81fb;
  wire al_e44d618;
  wire al_6ab58fb5;
  wire al_37c809df;
  wire al_1d552e04;
  wire al_307af410;
  wire al_1e561c50;
  wire al_9b855829;
  wire al_41381f51;
  wire al_2e700a59;
  wire al_e7a9a14d;
  wire al_6cdf2816;
  wire al_3370be13;
  wire al_c1d58f9c;
  wire al_7557c0dc;
  wire al_994b00c4;
  wire al_a783ebfd;
  wire al_51ab8bb8;
  wire al_1ed21a96;
  wire al_2c7a1247;
  wire al_fe00f314;
  wire al_db3c8a2c;
  wire al_4f9f38e2;
  wire al_4f1a9685;
  wire al_cca5b6a5;
  wire al_823fecd4;
  wire al_ccf401cd;
  wire al_735aa681;
  wire al_1180f8c0;
  wire al_a0088870;
  wire al_18337cf7;
  wire al_99f08586;
  wire al_bba5a10a;
  wire al_70b7c327;
  wire al_be034ab5;
  wire al_f205e138;
  wire al_d86c9f70;
  wire al_618737cb;
  wire al_f0947bb5;
  wire al_4290d1b8;
  wire al_8996909b;
  wire al_e1409b5e;
  wire al_2787c2b9;
  wire al_4cf5bca0;
  wire al_a396e89f;
  wire al_890eb5a1;
  wire al_63101725;
  wire al_949a133d;
  wire al_cc14f446;
  wire al_27161c58;
  wire al_e4f71d03;
  wire al_34aaf187;
  wire al_87b441ee;
  wire al_6ec43dd2;
  wire al_59c37d06;
  wire al_f7483e6d;
  wire al_1ff7640d;
  wire al_1c08f670;
  wire al_68c341e7;
  wire al_27717189;
  wire al_e3955cca;
  wire al_baa47a85;
  wire al_bffbe171;
  wire al_342f6170;
  wire al_dacef8ff;
  wire al_15c18023;
  wire al_8999d24b;
  wire al_3a7c57e3;
  wire al_bb167cdd;
  wire al_fe465555;
  wire al_76ee0125;
  wire al_aeadc72a;
  wire al_3e13fa86;
  wire al_1629ae4d;
  wire al_31732ee5;
  wire al_e3b877ad;
  wire al_1af0ad5e;
  wire al_e1d5aa87;
  wire al_a1ace55b;
  wire al_fa54303d;
  wire al_8aec7267;
  wire al_75c3c1c0;
  wire al_c8fffdaf;
  wire al_8769457b;
  wire al_1c648f36;
  wire al_af3abf3a;
  wire al_473186ca;
  wire al_33991d35;
  wire al_506bb8a;
  wire al_1973de82;
  wire al_1bae0f4e;
  wire al_7f95b06f;
  wire al_83c2aae7;
  wire al_1adec7e7;
  wire al_3714f7a3;
  wire al_23cb1fcc;
  wire al_407365eb;
  wire al_bcf9a5e2;
  wire al_4529840c;
  wire al_6333de40;
  wire al_d8bfe065;
  wire al_164531d8;
  wire al_20c70ab1;
  wire al_458cb894;
  wire al_88b7c5fc;
  wire al_8cf1eeca;
  wire al_6a75b886;
  wire al_c5c11e98;
  wire al_aa43251;
  wire al_db02221b;
  wire al_1217cf69;
  wire al_fdcd79c7;
  wire al_f50bd9c;
  wire al_2ef0a421;
  wire al_d9ec2230;
  wire al_49c3c8c7;
  wire al_40258be6;
  wire al_fc6a7e7a;
  wire al_755e05f8;
  wire al_604d05a2;
  wire al_53de47ce;
  wire al_fc5f2d2a;
  wire al_88f7ad44;
  wire al_d407324e;
  wire al_afc1b64;
  wire al_76e54a1a;
  wire al_aa509190;
  wire al_f766fdfa;
  wire al_379b9322;
  wire al_4df60ad5;
  wire al_8e2f2cc5;
  wire al_e2923d0b;
  wire al_5607a442;
  wire al_482a08f7;
  wire al_b3908a65;
  wire al_86d0105a;
  wire al_1c8c2124;
  wire al_adafc833;
  wire al_fb0d0f97;
  wire al_7fbfd2c7;
  wire al_63bd33e6;
  wire al_4c800f86;
  wire al_1b903e6a;
  wire al_35f01e82;
  wire al_fd6c10a8;
  wire al_fd9c8287;
  wire al_8587a543;
  wire al_6b181c0;
  wire al_90591ccb;
  wire al_5bf34257;
  wire al_43c0413c;
  wire al_d94de5f0;
  wire al_8f504dd9;
  wire al_7bf90fef;
  wire al_82626899;
  wire al_ec8f4956;
  wire al_d7d4dbcb;
  wire al_a97b8529;
  wire al_dc2d168e;
  wire al_8127333f;
  wire al_6dcc3ceb;
  wire al_495ff86c;
  wire al_7a7f52dd;
  wire al_a29e073;
  wire al_711bc49b;
  wire al_b256aea1;
  wire al_452179e4;
  wire al_64bdbb03;
  wire al_ec6037b6;
  wire al_8e038ddf;
  wire al_337e2949;
  wire al_84914f7c;
  wire al_99b7d851;
  wire al_b945c2ed;
  wire al_ccb46709;
  wire al_f1c0edfa;
  wire al_1e5502f4;
  wire al_2c28807a;
  wire al_153ccbd8;
  wire al_eae41b9d;
  wire al_45b5d05e;
  wire al_9f0f27fb;
  wire al_9e512d7f;
  wire al_d889aa1d;
  wire al_f751b948;
  wire al_37d9882e;
  wire al_7e094735;
  wire al_36697857;
  wire al_f817c39d;
  wire al_1041edd0;
  wire al_1a3cae1d;
  wire al_60cada77;
  wire al_97f75483;
  wire al_df62d485;
  wire al_19219cae;
  wire al_31650bb3;
  wire al_986ad8e6;
  wire al_d0cbf8c4;
  wire al_a4119c94;
  wire al_1ca6a854;
  wire al_d439eb63;
  wire al_e7647890;
  wire al_624c8b6f;
  wire al_a9406400;
  wire al_dbd330f5;
  wire al_5d31465b;
  wire al_c3d9ce92;
  wire al_1b655917;
  wire al_291f5813;
  wire al_35a8bfef;
  wire al_ad19785e;
  wire al_1c908f3d;
  wire al_fc6dfd0c;
  wire al_2e19f5ba;
  wire al_57e16e6f;
  wire al_d5f82e51;
  wire al_3fec348f;
  wire al_1ce50ae3;
  wire al_bf676c3e;
  wire al_a584e1fd;
  wire al_2086b792;
  wire al_1d703c48;
  wire al_d016a646;
  wire al_d376e8f0;
  wire al_e25f50ab;
  wire al_9befeaf3;
  wire al_6dd1a6b;
  wire al_ca75b795;
  wire al_2dc26b59;
  wire al_314de0e;
  wire al_84d6d5e6;
  wire al_70a55548;
  wire al_a51b1b3a;
  wire al_acb683b9;
  wire al_7f071305;
  wire al_a511ca2d;
  wire al_60c51ee3;
  wire al_c53dc261;
  wire al_e7834cb3;
  wire al_144281a5;
  wire al_dcaf20fc;
  wire al_ad53d9d0;
  wire al_ffec892d;
  wire al_d24d858b;
  wire al_6400d4de;
  wire al_e8e15f03;
  wire al_2014d3d9;
  wire al_39855db7;
  wire al_6230936a;
  wire al_aacd2311;
  wire al_c1b912e;
  wire al_48bec3d3;
  wire al_751a5b13;
  wire al_572dc31a;
  wire al_3b935332;
  wire al_c68dfd58;
  wire al_4e8c0a64;
  wire al_6a1aebd1;
  wire al_c9bfee53;
  wire al_7968b2a5;
  wire al_7c711acd;
  wire al_14e5d384;
  wire al_c6d1dc18;
  wire al_2b48f483;
  wire al_841146bf;
  wire al_3cbc9279;
  wire al_f3e1aff9;
  wire al_10307540;
  wire al_332cacdd;
  wire al_bfa502a9;
  wire al_a53ff9fc;
  wire al_8f82c712;
  wire al_82faa065;
  wire al_b7164eee;
  wire al_e3838f69;
  wire al_4965e5fa;
  wire al_71f17e1a;
  wire al_41ffdcd4;
  wire al_7afe69f4;
  wire al_74a15ab1;
  wire al_5ec57682;
  wire al_2da9429f;
  wire al_64bc3920;
  wire al_b39aa369;
  wire al_60993b86;
  wire al_edca2c86;
  wire al_711d3f5;
  wire al_3c3908e6;
  wire al_da959817;
  wire al_ef45b73e;
  wire al_f7e49aaa;
  wire al_f5bbf69e;
  wire al_a8b162ca;
  wire al_f474e268;
  wire al_8952b398;
  wire al_78512832;
  wire al_715827e7;
  wire al_740a6bb3;
  wire al_b17db8f;
  wire al_b1b43431;
  wire al_8e2b6222;
  wire al_7fea7bf;
  wire al_ff09d078;
  wire al_38f26a35;
  wire al_62d97d99;
  wire al_cf696ef0;
  wire al_ad22e376;
  wire al_a9336f5;
  wire al_30b5e311;
  wire al_2110386e;
  wire al_536b4576;
  wire al_3edda74b;
  wire al_dbe2baa6;
  wire al_8f15a934;
  wire al_b5e36a9;
  wire al_d976dda9;
  wire al_4596a396;
  wire al_59a83809;
  wire al_1bc55ab2;
  wire al_1c6db97d;
  wire al_68a14bd2;
  wire al_56997d45;
  wire al_982b355d;
  wire al_f16b3d6d;
  wire al_49c7fc0e;
  wire al_113d1401;
  wire al_8e145e50;
  wire al_4efdb29f;
  wire al_3e178366;
  wire al_56b3d928;
  wire al_66d47dbf;
  wire al_dc21b291;
  wire al_db67c2f5;
  wire al_e4f9c44c;
  wire al_d23bd93a;
  wire al_f7638b94;
  wire al_dc8505e1;
  wire al_134c8dab;
  wire al_78991444;
  wire al_ce826c89;
  wire al_175588ec;
  wire al_6aaeddf4;
  wire al_1430ac7c;
  wire al_9b5719ae;
  wire al_f2d1cf9;
  wire al_7be18307;
  wire al_8ab6e600;
  wire al_4974667d;
  wire al_fd84e521;
  wire al_1f5e6438;
  wire al_e410470b;
  wire al_587ea99f;
  wire al_6bff803e;
  wire al_2a3de543;
  wire al_5716efe6;
  wire al_70d272c9;
  wire al_7b32ad34;
  wire al_ab134353;
  wire al_3eaa9cdd;
  wire al_53669626;
  wire al_f452d0ae;
  wire al_edebc70b;
  wire al_e6700530;
  wire al_8d4887c7;
  wire al_aaacabd5;
  wire al_1ec4cd29;
  wire al_88a2bdf0;
  wire al_468d7712;
  wire al_1b37ba12;
  wire al_9c1262a5;
  wire al_fcec21f3;
  wire al_39bb30c0;
  wire al_d6e69fcf;
  wire al_3b01668f;
  wire al_1e78f688;
  wire al_13600bf4;
  wire al_5bb5921;
  wire al_a024e6ee;
  wire al_33c6f6;
  wire al_f9f3df5f;
  wire al_ebd95b94;
  wire al_522428e2;
  wire al_4690bf2e;
  wire al_f23520ad;
  wire al_d48745aa;
  wire al_a8508f7c;
  wire al_a50e12e0;
  wire al_221dcd70;
  wire al_1af55219;
  wire al_88de809d;
  wire al_d3c8ca1c;
  wire al_c39b1824;
  wire al_b89e105d;
  wire al_a2d9d6a;
  wire al_a0e3e4ed;
  wire al_215b7b3d;
  wire al_8d6efaba;
  wire al_114295f1;
  wire al_8e55a7af;
  wire al_9d9dbb20;
  wire al_6ab23518;
  wire al_968fd17c;
  wire al_4f2f7ae3;
  wire al_904a5dce;
  wire al_fc8b055a;

  assign gmii_tx_en = al_1a7bad30;
  assign gmii_tx_er = al_e5091a32;
  assign gmii_txd[7] = al_bb772f98[7];
  assign gmii_txd[6] = al_bb772f98[6];
  assign gmii_txd[5] = al_bb772f98[5];
  assign gmii_txd[4] = al_bb772f98[4];
  assign gmii_txd[3] = al_bb772f98[3];
  assign gmii_txd[2] = al_bb772f98[2];
  assign gmii_txd[1] = al_bb772f98[1];
  assign gmii_txd[0] = al_bb772f98[0];
  assign s_axi_awready = s_axi_wready;
  assign s_axi_bresp[1] = 1'b0;
  assign s_axi_bresp[0] = 1'b0;
  assign s_axi_rresp[1] = 1'b0;
  assign s_axi_rresp[0] = 1'b0;
  AL_DFF_X al_2f20b443 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_dad1457e),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(tx_status_vector[3]));
  AL_DFF_X al_6c7765cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f7d4c035),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_2bb2d81d));
  AL_DFF_X al_b270513d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5374577),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_678e4333));
  AL_MAP_LUT6 #(
    .EQN("(~F*E*~D*C*B*A)"),
    .INIT(64'h0000000000800000))
    al_44c81e3b (
    .a(al_4f0de751),
    .b(al_ba2c5d76),
    .c(rx_clk_en),
    .d(al_bd4c52f0[0]),
    .e(al_bd4c52f0[3]),
    .f(al_bd4c52f0[4]),
    .o(al_1a6b1e5a));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~((E*~D*~C*B))*~(F)+~(A)*(E*~D*~C*B)*~(F)+A*~((E*~D*~C*B))*F+~(A)*(E*~D*~C*B)*F+A*(E*~D*~C*B)*F)"),
    .INIT(64'haaaeaaaa55555555))
    al_20475d1a (
    .a(al_bd4c52f0[0]),
    .b(al_bd4c52f0[1]),
    .c(al_bd4c52f0[2]),
    .d(al_bd4c52f0[3]),
    .e(al_bd4c52f0[4]),
    .f(al_8b7d9749),
    .o(al_71becb96));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_41604787 (
    .a(al_71becb96),
    .b(al_4f0de751),
    .o(al_d002eac[0]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C@(D*B)))"),
    .INIT(16'h28a0))
    al_b765bf2a (
    .a(al_4f0de751),
    .b(al_bd4c52f0[0]),
    .c(al_bd4c52f0[1]),
    .d(al_8b7d9749),
    .o(al_d002eac[1]));
  AL_MAP_LUT5 #(
    .EQN("(A*(D@(E*C*B)))"),
    .INIT(32'h2a80aa00))
    al_b2adbb47 (
    .a(al_4f0de751),
    .b(al_bd4c52f0[0]),
    .c(al_bd4c52f0[1]),
    .d(al_bd4c52f0[2]),
    .e(al_8b7d9749),
    .o(al_d002eac[2]));
  AL_MAP_LUT5 #(
    .EQN("(A*(D@(E*C*B)))"),
    .INIT(32'h2a80aa00))
    al_92ca88d3 (
    .a(al_4f0de751),
    .b(al_ba2c5d76),
    .c(al_bd4c52f0[0]),
    .d(al_bd4c52f0[3]),
    .e(al_8b7d9749),
    .o(al_d002eac[3]));
  AL_MAP_LUT6 #(
    .EQN("(A*(E@(F*D*C*B)))"),
    .INIT(64'h2aaa8000aaaa0000))
    al_df16d585 (
    .a(al_4f0de751),
    .b(al_ba2c5d76),
    .c(al_bd4c52f0[0]),
    .d(al_bd4c52f0[3]),
    .e(al_bd4c52f0[4]),
    .f(al_8b7d9749),
    .o(al_d002eac[4]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_10b1f3b2 (
    .a(al_1feb4c09),
    .b(al_e2b7a540),
    .o(al_4f0de751));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_125bb27f (
    .a(al_14acaf34),
    .b(al_5160c8c2[1]),
    .c(al_5160c8c2[2]),
    .o(al_50f7b858));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~(B*A)))"),
    .INIT(16'hf080))
    al_31c96e92 (
    .a(al_50f7b858),
    .b(al_dc85d54),
    .c(al_4f0de751),
    .d(al_678e4333),
    .o(al_5374577));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_5abdde44 (
    .a(al_bd4c52f0[1]),
    .b(al_bd4c52f0[2]),
    .o(al_ba2c5d76));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    al_2ed27013 (
    .a(al_ba2c5d76),
    .b(al_bd4c52f0[0]),
    .c(al_bd4c52f0[3]),
    .d(al_bd4c52f0[4]),
    .o(al_dc85d54));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_8553d2a3 (
    .a(al_e8c856c9[4]),
    .b(al_e8c856c9[5]),
    .c(al_e8c856c9[6]),
    .d(al_e8c856c9[7]),
    .o(al_a700dfa6));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*A)"),
    .INIT(64'h0000000000000002))
    al_1d759451 (
    .a(al_5160c8c2[0]),
    .b(al_5160c8c2[3]),
    .c(al_5160c8c2[4]),
    .d(al_5160c8c2[5]),
    .e(al_5160c8c2[6]),
    .f(al_5160c8c2[7]),
    .o(al_74b73e47));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*B*A)"),
    .INIT(64'h0000000000000008))
    al_d5031047 (
    .a(al_74b73e47),
    .b(al_a700dfa6),
    .c(al_e8c856c9[0]),
    .d(al_e8c856c9[1]),
    .e(al_e8c856c9[2]),
    .f(al_e8c856c9[3]),
    .o(al_14acaf34));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    al_5eb082a2 (
    .a(al_7b7a3c37),
    .b(al_4f0de751),
    .c(al_2c28b3bd[0]),
    .d(al_5160c8c2[0]),
    .o(al_b9f27169[0]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    al_9087e751 (
    .a(al_d61cd20b),
    .b(al_4f0de751),
    .c(al_2c28b3bd[10]),
    .d(al_5160c8c2[2]),
    .o(al_b9f27169[10]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    al_71264a1e (
    .a(al_d61cd20b),
    .b(al_4f0de751),
    .c(al_2c28b3bd[11]),
    .d(al_5160c8c2[3]),
    .o(al_b9f27169[11]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    al_412f6fb2 (
    .a(al_d61cd20b),
    .b(al_4f0de751),
    .c(al_2c28b3bd[12]),
    .d(al_5160c8c2[4]),
    .o(al_b9f27169[12]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    al_fb2eadcd (
    .a(al_d61cd20b),
    .b(al_4f0de751),
    .c(al_2c28b3bd[13]),
    .d(al_5160c8c2[5]),
    .o(al_b9f27169[13]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    al_3f122568 (
    .a(al_d61cd20b),
    .b(al_4f0de751),
    .c(al_2c28b3bd[14]),
    .d(al_5160c8c2[6]),
    .o(al_b9f27169[14]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    al_10658ce9 (
    .a(al_d61cd20b),
    .b(al_4f0de751),
    .c(al_2c28b3bd[15]),
    .d(al_5160c8c2[7]),
    .o(al_b9f27169[15]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    al_d76a4096 (
    .a(al_7b7a3c37),
    .b(al_4f0de751),
    .c(al_2c28b3bd[1]),
    .d(al_5160c8c2[1]),
    .o(al_b9f27169[1]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    al_352934bb (
    .a(al_7b7a3c37),
    .b(al_4f0de751),
    .c(al_2c28b3bd[2]),
    .d(al_5160c8c2[2]),
    .o(al_b9f27169[2]));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*~B*A)"),
    .INIT(32'h00020000))
    al_cefae771 (
    .a(al_bd4c52f0[0]),
    .b(al_bd4c52f0[1]),
    .c(al_bd4c52f0[2]),
    .d(al_bd4c52f0[3]),
    .e(al_bd4c52f0[4]),
    .o(al_7b7a3c37));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    al_919659ab (
    .a(al_7b7a3c37),
    .b(al_4f0de751),
    .c(al_2c28b3bd[3]),
    .d(al_5160c8c2[3]),
    .o(al_b9f27169[3]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    al_30d6b71 (
    .a(al_7b7a3c37),
    .b(al_4f0de751),
    .c(al_2c28b3bd[4]),
    .d(al_5160c8c2[4]),
    .o(al_b9f27169[4]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    al_6897e62c (
    .a(al_7b7a3c37),
    .b(al_4f0de751),
    .c(al_2c28b3bd[5]),
    .d(al_5160c8c2[5]),
    .o(al_b9f27169[5]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    al_861508ea (
    .a(al_7b7a3c37),
    .b(al_4f0de751),
    .c(al_2c28b3bd[6]),
    .d(al_5160c8c2[6]),
    .o(al_b9f27169[6]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    al_36a4034a (
    .a(al_7b7a3c37),
    .b(al_4f0de751),
    .c(al_2c28b3bd[7]),
    .d(al_5160c8c2[7]),
    .o(al_b9f27169[7]));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*~B*~A)"),
    .INIT(32'h00010000))
    al_10306764 (
    .a(al_bd4c52f0[0]),
    .b(al_bd4c52f0[1]),
    .c(al_bd4c52f0[2]),
    .d(al_bd4c52f0[3]),
    .e(al_bd4c52f0[4]),
    .o(al_d61cd20b));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    al_5740deb3 (
    .a(al_d61cd20b),
    .b(al_4f0de751),
    .c(al_2c28b3bd[8]),
    .d(al_5160c8c2[0]),
    .o(al_b9f27169[8]));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    al_88d99a5a (
    .a(al_d61cd20b),
    .b(al_4f0de751),
    .c(al_2c28b3bd[9]),
    .d(al_5160c8c2[1]),
    .o(al_b9f27169[9]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~(B*~A)))"),
    .INIT(16'hf040))
    al_6e3c1a56 (
    .a(al_50f7b858),
    .b(al_dc85d54),
    .c(al_4f0de751),
    .d(al_2bb2d81d),
    .o(al_f7d4c035));
  AL_DFF_X al_5c9ffeb5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b9f27169[0]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_2c28b3bd[0]));
  AL_DFF_X al_ce67489 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b9f27169[9]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_2c28b3bd[9]));
  AL_DFF_X al_58c802c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b9f27169[10]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_2c28b3bd[10]));
  AL_DFF_X al_da56e0a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b9f27169[11]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_2c28b3bd[11]));
  AL_DFF_X al_c1e58cd3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b9f27169[12]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_2c28b3bd[12]));
  AL_DFF_X al_d169d3be (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b9f27169[13]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_2c28b3bd[13]));
  AL_DFF_X al_61f06c28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b9f27169[14]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_2c28b3bd[14]));
  AL_DFF_X al_62eb3a7b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b9f27169[15]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_2c28b3bd[15]));
  AL_DFF_X al_16c37b54 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b9f27169[1]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_2c28b3bd[1]));
  AL_DFF_X al_1f00f9b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b9f27169[2]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_2c28b3bd[2]));
  AL_DFF_X al_f57b00c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b9f27169[3]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_2c28b3bd[3]));
  AL_DFF_X al_d377c341 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b9f27169[4]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_2c28b3bd[4]));
  AL_DFF_X al_e5b35c6a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b9f27169[5]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_2c28b3bd[5]));
  AL_DFF_X al_c3d147e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b9f27169[6]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_2c28b3bd[6]));
  AL_DFF_X al_1290ad58 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b9f27169[7]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_2c28b3bd[7]));
  AL_DFF_X al_61ffc201 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b9f27169[8]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_2c28b3bd[8]));
  AL_DFF_X al_cdcf185 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5160c8c2[0]),
    .en(al_1a6b1e5a),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_e8c856c9[0]));
  AL_DFF_X al_fbda843c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5160c8c2[1]),
    .en(al_1a6b1e5a),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_e8c856c9[1]));
  AL_DFF_X al_f2621fde (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5160c8c2[2]),
    .en(al_1a6b1e5a),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_e8c856c9[2]));
  AL_DFF_X al_65c11fbe (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5160c8c2[3]),
    .en(al_1a6b1e5a),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_e8c856c9[3]));
  AL_DFF_X al_8c7c204 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5160c8c2[4]),
    .en(al_1a6b1e5a),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_e8c856c9[4]));
  AL_DFF_X al_666dffe5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5160c8c2[5]),
    .en(al_1a6b1e5a),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_e8c856c9[5]));
  AL_DFF_X al_8c953167 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5160c8c2[6]),
    .en(al_1a6b1e5a),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_e8c856c9[6]));
  AL_DFF_X al_349ce4cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5160c8c2[7]),
    .en(al_1a6b1e5a),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_e8c856c9[7]));
  AL_DFF_X al_94e94a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_d002eac[0]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_bd4c52f0[0]));
  AL_DFF_X al_2ea42c5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_d002eac[1]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_bd4c52f0[1]));
  AL_DFF_X al_6f6c052e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_d002eac[2]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_bd4c52f0[2]));
  AL_DFF_X al_445d7aae (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_d002eac[3]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_bd4c52f0[3]));
  AL_DFF_X al_b0075a80 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_d002eac[4]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_bd4c52f0[4]));
  AL_MAP_LUT5 #(
    .EQN("~(~D*~(E*C*~B*A))"),
    .INIT(32'hff20ff00))
    al_b93afce8 (
    .a(al_abc98a52),
    .b(al_2bb2d81d),
    .c(al_1feb4c09),
    .d(al_e2b7a540),
    .e(al_8b780845),
    .o(al_e8fc825c));
  AL_DFF_X al_5241f804 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e8fc825c),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_error_frame));
  AL_DFF_X al_35cc110e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_8b7d9749),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_data_vld));
  AL_DFF_X al_3e9ff589 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_2e1a2363),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_abc98a52));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D*~B*A))"),
    .INIT(16'hd0f0))
    al_8fe2ef13 (
    .a(al_abc98a52),
    .b(al_2bb2d81d),
    .c(al_1feb4c09),
    .d(al_8b780845),
    .o(al_7c94b9c5));
  AL_DFF_X al_e90cf8c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_7c94b9c5),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_correct_frame));
  AL_DFF_X al_1b46f63 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1feb4c09),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_d5df3ac1));
  AL_DFF_X al_84169261 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_d5df3ac1),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_53bc66bd));
  AL_DFF_X al_373c107 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_53bc66bd),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_d30618ea));
  AL_DFF_X al_36eb4c38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_9c3c5741),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_59f1a9e9));
  AL_DFF_X al_72609d39 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_6de80447),
    .en(al_b2ee3fbb),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_ec74b2dd));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_a400fa3a (
    .a(rx_clk_en),
    .b(al_1feb4c09),
    .o(al_b2ee3fbb));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*~A)"),
    .INIT(8'hfe))
    al_e453f29e (
    .a(al_53bc66bd),
    .b(al_d30618ea),
    .c(al_d5df3ac1),
    .o(al_9c3c5741));
  AL_DFF_X al_475b49d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_2c28b3bd[0]),
    .en(al_b2ee3fbb),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_a6672453[0]));
  AL_DFF_X al_30f7117e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_2c28b3bd[9]),
    .en(al_b2ee3fbb),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_a6672453[9]));
  AL_DFF_X al_f24a52ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_2c28b3bd[10]),
    .en(al_b2ee3fbb),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_a6672453[10]));
  AL_DFF_X al_c8332e2e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_2c28b3bd[11]),
    .en(al_b2ee3fbb),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_a6672453[11]));
  AL_DFF_X al_bd2b6d05 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_2c28b3bd[12]),
    .en(al_b2ee3fbb),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_a6672453[12]));
  AL_DFF_X al_ab1d15a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_2c28b3bd[13]),
    .en(al_b2ee3fbb),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_a6672453[13]));
  AL_DFF_X al_1c2b9e57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_2c28b3bd[14]),
    .en(al_b2ee3fbb),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_a6672453[14]));
  AL_DFF_X al_19012e36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_2c28b3bd[15]),
    .en(al_b2ee3fbb),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_a6672453[15]));
  AL_DFF_X al_af6f34e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_2c28b3bd[1]),
    .en(al_b2ee3fbb),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_a6672453[1]));
  AL_DFF_X al_1ce136d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_2c28b3bd[2]),
    .en(al_b2ee3fbb),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_a6672453[2]));
  AL_DFF_X al_bbdf49a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_2c28b3bd[3]),
    .en(al_b2ee3fbb),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_a6672453[3]));
  AL_DFF_X al_f81e09fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_2c28b3bd[4]),
    .en(al_b2ee3fbb),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_a6672453[4]));
  AL_DFF_X al_e62d1f2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_2c28b3bd[5]),
    .en(al_b2ee3fbb),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_a6672453[5]));
  AL_DFF_X al_5345a5e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_2c28b3bd[6]),
    .en(al_b2ee3fbb),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_a6672453[6]));
  AL_DFF_X al_13915ebd (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_2c28b3bd[7]),
    .en(al_b2ee3fbb),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_a6672453[7]));
  AL_DFF_X al_76994b4f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_2c28b3bd[8]),
    .en(al_b2ee3fbb),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_a6672453[8]));
  AL_DFF_X al_75d5369f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_fa26b745),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_6e8a0941));
  AL_DFF_X al_54aeeda9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_32868173),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_77b8d1cd));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_343e1d55 (
    .a(tx_data_en),
    .b(al_77b8d1cd),
    .o(tx_rdy));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    al_b108bf76 (
    .a(al_24ac8493[0]),
    .b(al_24ac8493[1]),
    .c(al_24ac8493[2]),
    .d(al_eb5c4882),
    .o(al_fa26b745));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(~B*~(~E*C*A)))"),
    .INIT(32'h00cc00ec))
    al_baf7af63 (
    .a(al_fa26b745),
    .b(tx_rdy),
    .c(tx_clk_en),
    .d(al_6b4499fc),
    .e(al_b984f6c1),
    .o(al_32868173));
  AL_DFF_X al_822c34ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5f71b9c1),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_bc147132));
  AL_DFF_X al_b10b45ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_data_en),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_ee74aec5));
  AL_DFF_X al_f003aeb7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c078e47f),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_20c861d8));
  AL_DFF_X al_14f65a23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_269c8a2f),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_77ced363));
  AL_DFF_X al_31d7dfb8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_80471da6),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_b984f6c1));
  AL_DFF_X al_e16b3019 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_6702ffbf),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_bc58b1b4));
  AL_MAP_LUT6 #(
    .EQN("(~B*~(A*~(F*~E*D)))"),
    .INIT(64'h1111331111111111))
    al_babc2e13 (
    .a(al_ee74aec5),
    .b(al_b984f6c1),
    .c(al_bc147132),
    .d(al_12358921),
    .e(al_68ba43d4),
    .f(al_9a8c459a),
    .o(al_c3d753a2));
  AL_MAP_LUT6 #(
    .EQN("(C*~B*~A*~(F*E*~D))"),
    .INIT(64'h1000101010101010))
    al_44d5d5ae (
    .a(al_c3d753a2),
    .b(al_d97145b1[1]),
    .c(al_d97145b1[2]),
    .d(al_1dee2dce[0]),
    .e(al_1dee2dce[1]),
    .f(al_1dee2dce[4]),
    .o(al_54e389b6));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(~A*~(E*~D*C)))"),
    .INIT(32'h22322222))
    al_97c273bf (
    .a(al_54e389b6),
    .b(al_d97145b1[0]),
    .c(al_d97145b1[1]),
    .d(al_d97145b1[2]),
    .e(al_6e8a0941),
    .o(al_2bf5454d));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(~E*~C*B*~A))"),
    .INIT(32'h00ff00fb))
    al_f82cb2fc (
    .a(al_20c861d8),
    .b(al_ee74aec5),
    .c(al_b984f6c1),
    .d(al_bc58b1b4),
    .e(al_89a3ef5a),
    .o(al_3956f95a));
  AL_MAP_LUT5 #(
    .EQN("(~D*(~(A)*B*~(C)*~(E)+~(A)*~(B)*C*~(E)+A*~(B)*C*~(E)+~(A)*B*~(C)*E))"),
    .INIT(32'h00040034))
    al_1c8d0fd2 (
    .a(al_3956f95a),
    .b(al_d97145b1[0]),
    .c(al_d97145b1[1]),
    .d(al_d97145b1[2]),
    .e(al_6e8a0941),
    .o(al_98b546cc));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hf5f5f0c5))
    al_faa77eaf (
    .a(al_54e389b6),
    .b(al_3956f95a),
    .c(al_d97145b1[0]),
    .d(al_d97145b1[1]),
    .e(al_d97145b1[2]),
    .o(al_8b27d348));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_7a67b387 (
    .a(tx_clk_en),
    .b(al_d97145b1[0]),
    .c(al_bc58b1b4),
    .o(al_92a04064));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_9739056 (
    .a(pause_req),
    .b(tx_clk_en),
    .o(al_f6b6167));
  AL_MAP_LUT4 #(
    .EQN("~(D*~C*B*A)"),
    .INIT(16'hf7ff))
    al_3cbbc7f1 (
    .a(al_2337d80f),
    .b(al_12358921),
    .c(al_68ba43d4),
    .d(al_9a8c459a),
    .o(al_269c8a2f));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~(B*A))"),
    .INIT(16'h0070))
    al_ff126423 (
    .a(al_20c861d8),
    .b(al_ee74aec5),
    .c(al_d97145b1[0]),
    .d(al_bc58b1b4),
    .o(al_dbdc14b4));
  AL_MAP_LUT6 #(
    .EQN("(E*~(A*~(F*~D*~C*B)))"),
    .INIT(64'h555d000055550000))
    al_375c42a9 (
    .a(al_dbdc14b4),
    .b(al_d97145b1[0]),
    .c(al_d97145b1[1]),
    .d(al_d97145b1[2]),
    .e(al_b984f6c1),
    .f(al_bc3d033e),
    .o(al_f4dbb19c));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~A*~(~(~E*~D)*~(C*B)))"),
    .INIT(64'hffffffffbfbfbfaa))
    al_9ad4af1f (
    .a(al_f4dbb19c),
    .b(al_269c8a2f),
    .c(al_ee74aec5),
    .d(al_bc58b1b4),
    .e(al_bc3d033e),
    .f(al_89a3ef5a),
    .o(al_80471da6));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*A))"),
    .INIT(8'hd0))
    al_a28fe597 (
    .a(al_269c8a2f),
    .b(al_20c861d8),
    .c(al_ee74aec5),
    .o(al_c078e47f));
  AL_MAP_LUT6 #(
    .EQN("(~(F*E*~D)*~(~C*~(B*A)))"),
    .INIT(64'hf800f8f8f8f8f8f8))
    al_8745b288 (
    .a(pause_req),
    .b(al_fc3c716f),
    .c(al_bc58b1b4),
    .d(al_1dee2dce[0]),
    .e(al_1dee2dce[1]),
    .f(al_1dee2dce[4]),
    .o(al_6702ffbf));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'h3a))
    al_e7d72cb5 (
    .a(al_21291e01),
    .b(al_bc58b1b4),
    .c(al_1dee2dce[0]),
    .o(al_7c53cb60[0]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h3ba0))
    al_7621f544 (
    .a(al_21291e01),
    .b(al_bc58b1b4),
    .c(al_1dee2dce[0]),
    .d(al_1dee2dce[1]),
    .o(al_7c53cb60[1]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B)*(D*C)*~(E)+A*B*(D*C)*~(E)+~(A)*~(B)*~((D*C))*E+A*~(B)*~((D*C))*E+A*B*~((D*C))*E+~(A)*~(B)*(D*C)*E+A*~(B)*(D*C)*E)"),
    .INIT(32'h3bbba000))
    al_e02d90ac (
    .a(al_21291e01),
    .b(al_bc58b1b4),
    .c(al_1dee2dce[0]),
    .d(al_1dee2dce[1]),
    .e(al_1dee2dce[2]),
    .o(al_7c53cb60[2]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*(E*D*C)*~(F)+A*B*(E*D*C)*~(F)+~(A)*~(B)*~((E*D*C))*F+A*~(B)*~((E*D*C))*F+A*B*~((E*D*C))*F+~(A)*~(B)*(E*D*C)*F+A*~(B)*(E*D*C)*F)"),
    .INIT(64'h3bbbbbbba0000000))
    al_79291c08 (
    .a(al_21291e01),
    .b(al_bc58b1b4),
    .c(al_1dee2dce[0]),
    .d(al_1dee2dce[1]),
    .e(al_1dee2dce[2]),
    .f(al_1dee2dce[3]),
    .o(al_7c53cb60[3]));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*B*A)"),
    .INIT(32'h00080000))
    al_d9ff8c1a (
    .a(al_1dee2dce[0]),
    .b(al_1dee2dce[1]),
    .c(al_1dee2dce[2]),
    .d(al_1dee2dce[3]),
    .e(al_1dee2dce[4]),
    .o(al_25ad8958));
  AL_MAP_LUT5 #(
    .EQN("(E*C*~A*~(~D*~B))"),
    .INIT(32'h50400000))
    al_81c4c8df (
    .a(al_25ad8958),
    .b(al_d97145b1[2]),
    .c(al_b984f6c1),
    .d(al_6e8a0941),
    .e(al_bc58b1b4),
    .o(al_21291e01));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_c57ee9a7 (
    .a(al_1dee2dce[0]),
    .b(al_1dee2dce[1]),
    .c(al_1dee2dce[2]),
    .d(al_1dee2dce[3]),
    .o(al_574485a3));
  AL_MAP_LUT4 #(
    .EQN("(A*B*~(C)*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D)"),
    .INIT(16'h2f88))
    al_76339080 (
    .a(al_21291e01),
    .b(al_574485a3),
    .c(al_bc58b1b4),
    .d(al_1dee2dce[4]),
    .o(al_7c53cb60[4]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00f0f0ccccaaaa))
    al_533a36ce (
    .a(al_9fdb6cdc[16]),
    .b(al_9fdb6cdc[24]),
    .c(al_9fdb6cdc[32]),
    .d(al_9fdb6cdc[40]),
    .e(al_1dee2dce[0]),
    .f(al_1dee2dce[1]),
    .o(al_36ab2fb9));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_ef7b46ed (
    .a(al_9fdb6cdc[0]),
    .b(al_9fdb6cdc[8]),
    .c(al_1dee2dce[0]),
    .o(al_d4f64f24));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hf000aaaa33f0000f))
    al_c275f0f2 (
    .a(al_36ab2fb9),
    .b(al_d4f64f24),
    .c(al_1dee2dce[0]),
    .d(al_1dee2dce[1]),
    .e(al_1dee2dce[2]),
    .f(al_1dee2dce[3]),
    .o(al_14405a50));
  AL_MAP_LUT6 #(
    .EQN("~(~((D*~(C)*~(E)+D*C*~(E)+~(D)*C*E+D*C*E)*B)*~(~F*A))"),
    .INIT(64'hc0c0cc00eaeaeeaa))
    al_dadeda31 (
    .a(al_14405a50),
    .b(al_d293a382),
    .c(al_27d2fc1a[0]),
    .d(al_27d2fc1a[8]),
    .e(al_1dee2dce[0]),
    .f(al_1dee2dce[4]),
    .o(al_9c572362[0]));
  AL_MAP_LUT5 #(
    .EQN("(D*(~(A)*~(B)*~(C)*~(E)+A*~(B)*~(C)*~(E)+~(A)*B*~(C)*~(E)+A*B*~(C)*~(E)+A*~(B)*~(C)*E+A*B*~(C)*E+~(A)*B*C*E+A*B*C*E))"),
    .INIT(32'hca000f00))
    al_c06c9d33 (
    .a(al_9fdb6cdc[1]),
    .b(al_9fdb6cdc[9]),
    .c(al_1dee2dce[0]),
    .d(al_1dee2dce[1]),
    .e(al_1dee2dce[2]),
    .o(al_e61a7e67));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00f0f0ccccaaaa))
    al_91aad6e0 (
    .a(al_9fdb6cdc[17]),
    .b(al_9fdb6cdc[25]),
    .c(al_9fdb6cdc[33]),
    .d(al_9fdb6cdc[41]),
    .e(al_1dee2dce[0]),
    .f(al_1dee2dce[1]),
    .o(al_b47e09b3));
  AL_MAP_LUT5 #(
    .EQN("(~E*(B*~((~C*A))*~(D)+B*(~C*A)*~(D)+~(B)*(~C*A)*D+B*(~C*A)*D))"),
    .INIT(32'h00000acc))
    al_614f4aca (
    .a(al_b47e09b3),
    .b(al_e61a7e67),
    .c(al_1dee2dce[2]),
    .d(al_1dee2dce[3]),
    .e(al_1dee2dce[4]),
    .o(al_6219a09a));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(B*(D*~(C)*~(E)+D*C*~(E)+~(D)*C*E+D*C*E)))"),
    .INIT(32'heaeaeeaa))
    al_e93289bb (
    .a(al_6219a09a),
    .b(al_d293a382),
    .c(al_27d2fc1a[1]),
    .d(al_27d2fc1a[9]),
    .e(al_1dee2dce[0]),
    .o(al_9c572362[1]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00f0f0ccccaaaa))
    al_ea161fc2 (
    .a(al_9fdb6cdc[18]),
    .b(al_9fdb6cdc[26]),
    .c(al_9fdb6cdc[34]),
    .d(al_9fdb6cdc[42]),
    .e(al_1dee2dce[0]),
    .f(al_1dee2dce[1]),
    .o(al_91e39671));
  AL_MAP_LUT6 #(
    .EQN("(~((D*~(E)*~(F)+D*E*~(F)+~(D)*E*F+D*E*F)*B)*~(C*A))"),
    .INIT(64'h13135f5f135f135f))
    al_5534bfc9 (
    .a(al_91e39671),
    .b(al_57e58431),
    .c(al_776d5772),
    .d(al_9fdb6cdc[2]),
    .e(al_9fdb6cdc[10]),
    .f(al_1dee2dce[0]),
    .o(al_5f618b63));
  AL_MAP_LUT6 #(
    .EQN("~(~((D*~(C)*~(E)+D*C*~(E)+~(D)*C*E+D*C*E)*B)*~(~F*~A))"),
    .INIT(64'hc0c0cc00d5d5dd55))
    al_1520dff9 (
    .a(al_5f618b63),
    .b(al_d293a382),
    .c(al_27d2fc1a[2]),
    .d(al_27d2fc1a[10]),
    .e(al_1dee2dce[0]),
    .f(al_1dee2dce[4]),
    .o(al_9c572362[2]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00f0f0ccccaaaa))
    al_1e0ab436 (
    .a(al_9fdb6cdc[19]),
    .b(al_9fdb6cdc[27]),
    .c(al_9fdb6cdc[35]),
    .d(al_9fdb6cdc[43]),
    .e(al_1dee2dce[0]),
    .f(al_1dee2dce[1]),
    .o(al_88c8ee13));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_3a3554e1 (
    .a(al_9fdb6cdc[3]),
    .b(al_9fdb6cdc[11]),
    .c(al_1dee2dce[0]),
    .o(al_b8dbdfec));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hf0553fff))
    al_df38b273 (
    .a(al_88c8ee13),
    .b(al_b8dbdfec),
    .c(al_1dee2dce[1]),
    .d(al_1dee2dce[2]),
    .e(al_1dee2dce[3]),
    .o(al_988cc37d));
  AL_MAP_LUT6 #(
    .EQN("~(~((D*~(C)*~(E)+D*C*~(E)+~(D)*C*E+D*C*E)*B)*~(~F*~A))"),
    .INIT(64'hc0c0cc00d5d5dd55))
    al_9ab0a376 (
    .a(al_988cc37d),
    .b(al_d293a382),
    .c(al_27d2fc1a[3]),
    .d(al_27d2fc1a[11]),
    .e(al_1dee2dce[0]),
    .f(al_1dee2dce[4]),
    .o(al_9c572362[3]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00f0f0ccccaaaa))
    al_718d91bd (
    .a(al_9fdb6cdc[20]),
    .b(al_9fdb6cdc[28]),
    .c(al_9fdb6cdc[36]),
    .d(al_9fdb6cdc[44]),
    .e(al_1dee2dce[0]),
    .f(al_1dee2dce[1]),
    .o(al_7bcff3b9));
  AL_MAP_LUT6 #(
    .EQN("(~((D*~(E)*~(F)+D*E*~(F)+~(D)*E*F+D*E*F)*B)*~(C*A))"),
    .INIT(64'h13135f5f135f135f))
    al_15527831 (
    .a(al_7bcff3b9),
    .b(al_57e58431),
    .c(al_776d5772),
    .d(al_9fdb6cdc[4]),
    .e(al_9fdb6cdc[12]),
    .f(al_1dee2dce[0]),
    .o(al_4bb8f8b3));
  AL_MAP_LUT6 #(
    .EQN("~(~((D*~(C)*~(E)+D*C*~(E)+~(D)*C*E+D*C*E)*B)*~(~F*~A))"),
    .INIT(64'hc0c0cc00d5d5dd55))
    al_8ea0220c (
    .a(al_4bb8f8b3),
    .b(al_d293a382),
    .c(al_27d2fc1a[4]),
    .d(al_27d2fc1a[12]),
    .e(al_1dee2dce[0]),
    .f(al_1dee2dce[4]),
    .o(al_9c572362[4]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_b06a7f32 (
    .a(al_1dee2dce[1]),
    .b(al_1dee2dce[2]),
    .c(al_1dee2dce[3]),
    .o(al_57e58431));
  AL_MAP_LUT6 #(
    .EQN("~(~((D*~(C)*~(E)+D*C*~(E)+~(D)*C*E+D*C*E)*B)*~(~F*~A))"),
    .INIT(64'hc0c0cc00d5d5dd55))
    al_6520cc92 (
    .a(al_be08372),
    .b(al_d293a382),
    .c(al_27d2fc1a[5]),
    .d(al_27d2fc1a[13]),
    .e(al_1dee2dce[0]),
    .f(al_1dee2dce[4]),
    .o(al_9c572362[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_ddf2ee8c (
    .a(al_1dee2dce[2]),
    .b(al_1dee2dce[3]),
    .o(al_776d5772));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    al_b42d5e15 (
    .a(al_1dee2dce[1]),
    .b(al_1dee2dce[2]),
    .c(al_1dee2dce[3]),
    .d(al_1dee2dce[4]),
    .o(al_d293a382));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00f0f0ccccaaaa))
    al_49dbb2e3 (
    .a(al_9fdb6cdc[21]),
    .b(al_9fdb6cdc[29]),
    .c(al_9fdb6cdc[37]),
    .d(al_9fdb6cdc[45]),
    .e(al_1dee2dce[0]),
    .f(al_1dee2dce[1]),
    .o(al_9d9cd237));
  AL_MAP_LUT6 #(
    .EQN("(~((D*~(E)*~(F)+D*E*~(F)+~(D)*E*F+D*E*F)*B)*~(C*A))"),
    .INIT(64'h13135f5f135f135f))
    al_cb36e1a6 (
    .a(al_9d9cd237),
    .b(al_57e58431),
    .c(al_776d5772),
    .d(al_9fdb6cdc[5]),
    .e(al_9fdb6cdc[13]),
    .f(al_1dee2dce[0]),
    .o(al_be08372));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h35f0))
    al_e0c89020 (
    .a(al_9fdb6cdc[6]),
    .b(al_9fdb6cdc[14]),
    .c(al_1dee2dce[0]),
    .d(al_1dee2dce[2]),
    .o(al_6f2ddcc1));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00f0f0ccccaaaa))
    al_27ae822 (
    .a(al_9fdb6cdc[22]),
    .b(al_9fdb6cdc[30]),
    .c(al_9fdb6cdc[38]),
    .d(al_9fdb6cdc[46]),
    .e(al_1dee2dce[0]),
    .f(al_1dee2dce[1]),
    .o(al_ed22e70c));
  AL_MAP_LUT5 #(
    .EQN("~((C*~B)*~((~D*A))*~(E)+(C*~B)*(~D*A)*~(E)+~((C*~B))*(~D*A)*E+(C*~B)*(~D*A)*E)"),
    .INIT(32'hff55cfcf))
    al_1b401a91 (
    .a(al_ed22e70c),
    .b(al_6f2ddcc1),
    .c(al_1dee2dce[1]),
    .d(al_1dee2dce[2]),
    .e(al_1dee2dce[3]),
    .o(al_cde2200a));
  AL_MAP_LUT6 #(
    .EQN("~(~((D*~(C)*~(E)+D*C*~(E)+~(D)*C*E+D*C*E)*B)*~(~F*~A))"),
    .INIT(64'hc0c0cc00d5d5dd55))
    al_4b441b6e (
    .a(al_cde2200a),
    .b(al_d293a382),
    .c(al_27d2fc1a[6]),
    .d(al_27d2fc1a[14]),
    .e(al_1dee2dce[0]),
    .f(al_1dee2dce[4]),
    .o(al_9c572362[6]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT(16'h88a0))
    al_70e2a55d (
    .a(al_d293a382),
    .b(al_27d2fc1a[7]),
    .c(al_27d2fc1a[15]),
    .d(al_1dee2dce[0]),
    .o(al_81b1fe1c));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00f0f0ccccaaaa))
    al_36a6897d (
    .a(al_9fdb6cdc[23]),
    .b(al_9fdb6cdc[31]),
    .c(al_9fdb6cdc[39]),
    .d(al_9fdb6cdc[47]),
    .e(al_1dee2dce[0]),
    .f(al_1dee2dce[1]),
    .o(al_83ef8a4e));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfff0ffff35fff00f))
    al_96ec504b (
    .a(al_9fdb6cdc[7]),
    .b(al_9fdb6cdc[15]),
    .c(al_1dee2dce[0]),
    .d(al_1dee2dce[1]),
    .e(al_1dee2dce[2]),
    .f(al_1dee2dce[3]),
    .o(al_bde4ed05));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(~E*~(C*~(D*B))))"),
    .INIT(32'haaaaefaf))
    al_7ad4f27a (
    .a(al_81b1fe1c),
    .b(al_83ef8a4e),
    .c(al_bde4ed05),
    .d(al_776d5772),
    .e(al_1dee2dce[4]),
    .o(al_9c572362[7]));
  AL_MAP_LUT6 #(
    .EQN("(~((~D*~C*~B))*~(E)*~((~F*~A))+(~D*~C*~B)*~(E)*~((~F*~A))+(~D*~C*~B)*E*~((~F*~A))+~((~D*~C*~B))*~(E)*(~F*~A)+(~D*~C*~B)*E*(~F*~A))"),
    .INIT(64'h0003ffff0003fffe))
    al_bb263305 (
    .a(al_1dee2dce[0]),
    .b(al_1dee2dce[1]),
    .c(al_1dee2dce[2]),
    .d(al_1dee2dce[3]),
    .e(al_1dee2dce[4]),
    .f(al_77ced363),
    .o(al_5f71b9c1));
  AL_DFF_X al_57367d97 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_8b27d348),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_d97145b1[0]));
  AL_DFF_X al_125ece25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_98b546cc),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_d97145b1[1]));
  AL_DFF_X al_90e811e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2bf5454d),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_d97145b1[2]));
  AL_DFF_X al_7581cb8f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_868a1cad[0]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[0]));
  AL_DFF_X al_2608eb21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_868a1cad[9]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[9]));
  AL_DFF_X al_f28cca76 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_868a1cad[10]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[10]));
  AL_DFF_X al_7e4da8fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_868a1cad[11]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[11]));
  AL_DFF_X al_eb3becc5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_868a1cad[12]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[12]));
  AL_DFF_X al_ca049f95 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_868a1cad[13]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[13]));
  AL_DFF_X al_791416fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_868a1cad[14]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[14]));
  AL_DFF_X al_cccbb35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_868a1cad[15]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[15]));
  AL_DFF_X al_9b0f747d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_868a1cad[16]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[16]));
  AL_DFF_X al_b98e2891 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_868a1cad[17]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[17]));
  AL_DFF_X al_3facc4e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_868a1cad[18]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[18]));
  AL_DFF_X al_3f13e4de (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_868a1cad[1]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[1]));
  AL_DFF_X al_e63a2edf (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_868a1cad[19]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[19]));
  AL_DFF_X al_56678233 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_868a1cad[20]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[20]));
  AL_DFF_X al_4fff4dc7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_868a1cad[21]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[21]));
  AL_DFF_X al_41bbe2e1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_868a1cad[22]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[22]));
  AL_DFF_X al_9965bf31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_868a1cad[23]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[23]));
  AL_DFF_X al_2b541ccb (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_868a1cad[24]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[24]));
  AL_DFF_X al_f15b9b9d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_868a1cad[25]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[25]));
  AL_DFF_X al_1357f4a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_868a1cad[26]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[26]));
  AL_DFF_X al_6c748ea2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_868a1cad[27]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[27]));
  AL_DFF_X al_ee3490fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_868a1cad[28]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[28]));
  AL_DFF_X al_e175076f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_868a1cad[2]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[2]));
  AL_DFF_X al_74768004 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_868a1cad[29]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[29]));
  AL_DFF_X al_62271c7e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_868a1cad[30]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[30]));
  AL_DFF_X al_fa329ace (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_868a1cad[31]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[31]));
  AL_DFF_X al_922a2537 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cd0aa0ee[0]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[32]));
  AL_DFF_X al_cfd7f589 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cd0aa0ee[1]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[33]));
  AL_DFF_X al_9e2e282 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cd0aa0ee[2]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[34]));
  AL_DFF_X al_3b9c411a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cd0aa0ee[3]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[35]));
  AL_DFF_X al_8989f43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cd0aa0ee[4]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[36]));
  AL_DFF_X al_20f4da30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cd0aa0ee[5]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[37]));
  AL_DFF_X al_4951beba (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cd0aa0ee[6]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[38]));
  AL_DFF_X al_3e9eb16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_868a1cad[3]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[3]));
  AL_DFF_X al_a8e0b69a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cd0aa0ee[7]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[39]));
  AL_DFF_X al_ac70782e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cd0aa0ee[8]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[40]));
  AL_DFF_X al_70b214f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cd0aa0ee[9]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[41]));
  AL_DFF_X al_6facc640 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cd0aa0ee[10]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[42]));
  AL_DFF_X al_d11be325 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cd0aa0ee[11]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[43]));
  AL_DFF_X al_8df2c165 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cd0aa0ee[12]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[44]));
  AL_DFF_X al_566a16b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cd0aa0ee[13]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[45]));
  AL_DFF_X al_46c80738 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cd0aa0ee[14]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[46]));
  AL_DFF_X al_f196c5ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cd0aa0ee[15]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[47]));
  AL_DFF_X al_b957fd10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_868a1cad[4]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[4]));
  AL_DFF_X al_6dfe5293 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_868a1cad[5]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[5]));
  AL_DFF_X al_e319034d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_868a1cad[6]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[6]));
  AL_DFF_X al_14968b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_868a1cad[7]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[7]));
  AL_DFF_X al_f306acd9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_868a1cad[8]),
    .en(al_92a04064),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9fdb6cdc[8]));
  AL_DFF_X al_36505cac (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(pause_val[0]),
    .en(al_f6b6167),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_27d2fc1a[0]));
  AL_DFF_X al_4dcb569a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(pause_val[9]),
    .en(al_f6b6167),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_27d2fc1a[9]));
  AL_DFF_X al_aebf3412 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(pause_val[10]),
    .en(al_f6b6167),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_27d2fc1a[10]));
  AL_DFF_X al_1fe440a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(pause_val[11]),
    .en(al_f6b6167),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_27d2fc1a[11]));
  AL_DFF_X al_d9bdf33 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(pause_val[12]),
    .en(al_f6b6167),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_27d2fc1a[12]));
  AL_DFF_X al_5a132143 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(pause_val[13]),
    .en(al_f6b6167),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_27d2fc1a[13]));
  AL_DFF_X al_f9fd80eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(pause_val[14]),
    .en(al_f6b6167),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_27d2fc1a[14]));
  AL_DFF_X al_b167955b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(pause_val[15]),
    .en(al_f6b6167),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_27d2fc1a[15]));
  AL_DFF_X al_260c3242 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(pause_val[1]),
    .en(al_f6b6167),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_27d2fc1a[1]));
  AL_DFF_X al_14467148 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(pause_val[2]),
    .en(al_f6b6167),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_27d2fc1a[2]));
  AL_DFF_X al_d617d35e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(pause_val[3]),
    .en(al_f6b6167),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_27d2fc1a[3]));
  AL_DFF_X al_15949f23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(pause_val[4]),
    .en(al_f6b6167),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_27d2fc1a[4]));
  AL_DFF_X al_2e7575b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(pause_val[5]),
    .en(al_f6b6167),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_27d2fc1a[5]));
  AL_DFF_X al_86400697 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(pause_val[6]),
    .en(al_f6b6167),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_27d2fc1a[6]));
  AL_DFF_X al_78d3ca9c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(pause_val[7]),
    .en(al_f6b6167),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_27d2fc1a[7]));
  AL_DFF_X al_8eb167b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(pause_val[8]),
    .en(al_f6b6167),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_27d2fc1a[8]));
  AL_DFF_X al_6c0c811c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_7c53cb60[0]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_1dee2dce[0]));
  AL_DFF_X al_b63a3ceb (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_7c53cb60[1]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_1dee2dce[1]));
  AL_DFF_X al_3ecc0937 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_7c53cb60[2]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_1dee2dce[2]));
  AL_DFF_X al_65acc8cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_7c53cb60[3]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_1dee2dce[3]));
  AL_DFF_X al_17bf3296 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_7c53cb60[4]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_1dee2dce[4]));
  AL_DFF_X al_cdcb5978 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9c572362[0]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_45ed4524[0]));
  AL_DFF_X al_fd4f7b90 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9c572362[1]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_45ed4524[1]));
  AL_DFF_X al_5c978bd1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9c572362[2]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_45ed4524[2]));
  AL_DFF_X al_28b4b361 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9c572362[3]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_45ed4524[3]));
  AL_DFF_X al_c37b4171 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9c572362[4]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_45ed4524[4]));
  AL_DFF_X al_9f501638 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9c572362[5]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_45ed4524[5]));
  AL_DFF_X al_a457a84e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9c572362[6]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_45ed4524[6]));
  AL_DFF_X al_a2f82364 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9c572362[7]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_45ed4524[7]));
  AL_DFF_X al_fc308f43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_206f470e),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(tx_collision));
  AL_DFF_X al_cbfae94b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_3fd53f68),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_fc3c716f));
  AL_DFF_X al_4717599 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_bc3d033e),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_adcb0cbd));
  AL_DFF_X al_86f15ce7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_27893604),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_bc3d033e));
  AL_DFF_X al_6a29f89b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_dd6bc6a),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_b1d5fd9b));
  AL_DFF_X al_4d2d7ed7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4e0a4dc5),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_89a3ef5a));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_6a0c3e6 (
    .a(al_a6672453[0]),
    .b(al_a6672453[1]),
    .c(al_a6672453[2]),
    .d(al_a6672453[3]),
    .o(al_c2dc89e9));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_de73911d (
    .a(al_a6672453[12]),
    .b(al_a6672453[13]),
    .c(al_a6672453[14]),
    .d(al_a6672453[15]),
    .o(al_7541e92c));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    al_7d74919b (
    .a(al_7541e92c),
    .b(al_a6672453[8]),
    .c(al_a6672453[9]),
    .d(al_a6672453[10]),
    .e(al_a6672453[11]),
    .o(al_6df60a04));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*B*A)"),
    .INIT(64'h0000000000000008))
    al_5724ae07 (
    .a(al_6df60a04),
    .b(al_c2dc89e9),
    .c(al_a6672453[4]),
    .d(al_a6672453[5]),
    .e(al_a6672453[6]),
    .f(al_a6672453[7]),
    .o(al_e98fadb));
  AL_MAP_LUT4 #(
    .EQN("~(~(~D*C)*~(A)*~(B)+~(~D*C)*A*~(B)+~(~(~D*C))*A*B+~(~D*C)*A*B)"),
    .INIT(16'h4474))
    al_68ed9cfe (
    .a(al_e98fadb),
    .b(al_62884f47),
    .c(al_bc3d033e),
    .d(al_89a3ef5a),
    .o(al_27893604));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_b3ff9ada (
    .a(al_ac3dcbf8[0]),
    .b(al_ac3dcbf8[3]),
    .c(al_ac3dcbf8[4]),
    .d(al_ac3dcbf8[5]),
    .e(al_ac3dcbf8[6]),
    .f(al_ac3dcbf8[7]),
    .o(al_d890a7e6));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_da894dde (
    .a(al_ac3dcbf8[8]),
    .b(al_ac3dcbf8[11]),
    .c(al_ac3dcbf8[12]),
    .d(al_ac3dcbf8[13]),
    .e(al_ac3dcbf8[14]),
    .f(al_ac3dcbf8[15]),
    .o(al_1ca8afe3));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*B*A)"),
    .INIT(64'h0000000000000008))
    al_80ee30c6 (
    .a(al_d890a7e6),
    .b(al_1ca8afe3),
    .c(al_ac3dcbf8[1]),
    .d(al_ac3dcbf8[2]),
    .e(al_ac3dcbf8[9]),
    .f(al_ac3dcbf8[10]),
    .o(al_8027e03));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*~(C*B)))"),
    .INIT(16'h5540))
    al_1bab4fb2 (
    .a(al_8027e03),
    .b(al_d97145b1[0]),
    .c(al_adcb0cbd),
    .d(al_89a3ef5a),
    .o(al_4e0a4dc5));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    al_8d154e7e (
    .a(al_d97145b1[0]),
    .b(al_bc3d033e),
    .c(al_38c57749[0]),
    .o(al_9868190b[0]));
  AL_MAP_LUT4 #(
    .EQN("((D@C)*~(B*A))"),
    .INIT(16'h0770))
    al_4526433f (
    .a(al_d97145b1[0]),
    .b(al_bc3d033e),
    .c(al_38c57749[0]),
    .d(al_38c57749[1]),
    .o(al_9868190b[1]));
  AL_MAP_LUT5 #(
    .EQN("((E@(D*C))*~(B*A))"),
    .INIT(32'h07777000))
    al_33684e82 (
    .a(al_d97145b1[0]),
    .b(al_bc3d033e),
    .c(al_38c57749[0]),
    .d(al_38c57749[1]),
    .e(al_38c57749[2]),
    .o(al_9868190b[2]));
  AL_MAP_LUT6 #(
    .EQN("((F@(E*D*C))*~(B*A))"),
    .INIT(64'h0777777770000000))
    al_2830d1f6 (
    .a(al_d97145b1[0]),
    .b(al_bc3d033e),
    .c(al_38c57749[0]),
    .d(al_38c57749[1]),
    .e(al_38c57749[2]),
    .f(al_38c57749[3]),
    .o(al_9868190b[3]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*(D@A))"),
    .INIT(16'h152a))
    al_40c6be1c (
    .a(al_633f8ef2),
    .b(al_d97145b1[0]),
    .c(al_bc3d033e),
    .d(al_38c57749[4]),
    .o(al_9868190b[4]));
  AL_MAP_LUT5 #(
    .EQN("(~(C*B)*(E@(D*A)))"),
    .INIT(32'h153f2a00))
    al_d9558488 (
    .a(al_633f8ef2),
    .b(al_d97145b1[0]),
    .c(al_bc3d033e),
    .d(al_38c57749[4]),
    .e(al_38c57749[5]),
    .o(al_9868190b[5]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_7520e0ba (
    .a(al_b746bad7),
    .b(al_62884f47),
    .c(al_a6672453[0]),
    .d(al_ac3dcbf8[0]),
    .e(al_dd86ad38[0]),
    .o(al_a128253b[0]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_25bc792d (
    .a(al_b746bad7),
    .b(al_62884f47),
    .c(al_a6672453[10]),
    .d(al_ac3dcbf8[10]),
    .e(al_dd86ad38[10]),
    .o(al_a128253b[10]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_2e0a1c44 (
    .a(al_b746bad7),
    .b(al_62884f47),
    .c(al_a6672453[11]),
    .d(al_ac3dcbf8[11]),
    .e(al_dd86ad38[11]),
    .o(al_a128253b[11]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_6e8ea480 (
    .a(al_b746bad7),
    .b(al_62884f47),
    .c(al_a6672453[12]),
    .d(al_ac3dcbf8[12]),
    .e(al_dd86ad38[12]),
    .o(al_a128253b[12]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_355a293f (
    .a(al_b746bad7),
    .b(al_62884f47),
    .c(al_a6672453[13]),
    .d(al_ac3dcbf8[13]),
    .e(al_dd86ad38[13]),
    .o(al_a128253b[13]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_177f343f (
    .a(al_38c57749[0]),
    .b(al_38c57749[1]),
    .c(al_38c57749[2]),
    .d(al_38c57749[3]),
    .o(al_633f8ef2));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    al_1834cbfd (
    .a(al_ec74b2dd),
    .b(al_b1d5fd9b),
    .c(al_dd6bc6a),
    .o(al_62884f47));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*C*~B*A)"),
    .INIT(32'h00200000))
    al_d0601ebc (
    .a(al_633f8ef2),
    .b(al_bc3d033e),
    .c(al_89a3ef5a),
    .d(al_38c57749[4]),
    .e(al_38c57749[5]),
    .o(al_b746bad7));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_7ad5e93 (
    .a(al_b746bad7),
    .b(al_62884f47),
    .c(al_a6672453[14]),
    .d(al_ac3dcbf8[14]),
    .e(al_dd86ad38[14]),
    .o(al_a128253b[14]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_c1caf22b (
    .a(al_b746bad7),
    .b(al_62884f47),
    .c(al_a6672453[15]),
    .d(al_ac3dcbf8[15]),
    .e(al_dd86ad38[15]),
    .o(al_a128253b[15]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_6bc63f89 (
    .a(al_b746bad7),
    .b(al_62884f47),
    .c(al_a6672453[1]),
    .d(al_ac3dcbf8[1]),
    .e(al_dd86ad38[1]),
    .o(al_a128253b[1]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_929a0054 (
    .a(al_b746bad7),
    .b(al_62884f47),
    .c(al_a6672453[2]),
    .d(al_ac3dcbf8[2]),
    .e(al_dd86ad38[2]),
    .o(al_a128253b[2]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_88032f2f (
    .a(al_b746bad7),
    .b(al_62884f47),
    .c(al_a6672453[3]),
    .d(al_ac3dcbf8[3]),
    .e(al_dd86ad38[3]),
    .o(al_a128253b[3]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_d60c9fb8 (
    .a(al_b746bad7),
    .b(al_62884f47),
    .c(al_a6672453[4]),
    .d(al_ac3dcbf8[4]),
    .e(al_dd86ad38[4]),
    .o(al_a128253b[4]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_6dcea23a (
    .a(al_b746bad7),
    .b(al_62884f47),
    .c(al_a6672453[5]),
    .d(al_ac3dcbf8[5]),
    .e(al_dd86ad38[5]),
    .o(al_a128253b[5]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_ff22a512 (
    .a(al_b746bad7),
    .b(al_62884f47),
    .c(al_a6672453[6]),
    .d(al_ac3dcbf8[6]),
    .e(al_dd86ad38[6]),
    .o(al_a128253b[6]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_3d62e7f7 (
    .a(al_b746bad7),
    .b(al_62884f47),
    .c(al_a6672453[7]),
    .d(al_ac3dcbf8[7]),
    .e(al_dd86ad38[7]),
    .o(al_a128253b[7]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_afef5244 (
    .a(al_b746bad7),
    .b(al_62884f47),
    .c(al_a6672453[8]),
    .d(al_ac3dcbf8[8]),
    .e(al_dd86ad38[8]),
    .o(al_a128253b[8]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_a4b14018 (
    .a(al_b746bad7),
    .b(al_62884f47),
    .c(al_a6672453[9]),
    .d(al_ac3dcbf8[9]),
    .e(al_dd86ad38[9]),
    .o(al_a128253b[9]));
  AL_DFF_X al_632d0da7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a128253b[0]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_ac3dcbf8[0]));
  AL_DFF_X al_7336bcf4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a128253b[9]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_ac3dcbf8[9]));
  AL_DFF_X al_ae070c3c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a128253b[10]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_ac3dcbf8[10]));
  AL_DFF_X al_88e3c458 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a128253b[11]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_ac3dcbf8[11]));
  AL_DFF_X al_639341ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a128253b[12]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_ac3dcbf8[12]));
  AL_DFF_X al_2345b94d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a128253b[13]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_ac3dcbf8[13]));
  AL_DFF_X al_85e2468d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a128253b[14]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_ac3dcbf8[14]));
  AL_DFF_X al_77577bd0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a128253b[15]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_ac3dcbf8[15]));
  AL_DFF_X al_5a8416f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a128253b[1]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_ac3dcbf8[1]));
  AL_DFF_X al_b58b0998 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a128253b[2]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_ac3dcbf8[2]));
  AL_DFF_X al_ab47471e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a128253b[3]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_ac3dcbf8[3]));
  AL_DFF_X al_3e326685 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a128253b[4]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_ac3dcbf8[4]));
  AL_DFF_X al_a55541a1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a128253b[5]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_ac3dcbf8[5]));
  AL_DFF_X al_3167bacf (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a128253b[6]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_ac3dcbf8[6]));
  AL_DFF_X al_5d19c132 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a128253b[7]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_ac3dcbf8[7]));
  AL_DFF_X al_fe8817d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a128253b[8]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_ac3dcbf8[8]));
  AL_DFF_X al_e430d3b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9868190b[0]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_38c57749[0]));
  AL_DFF_X al_93013923 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9868190b[1]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_38c57749[1]));
  AL_DFF_X al_1adbf48e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9868190b[2]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_38c57749[2]));
  AL_DFF_X al_a8251b34 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9868190b[3]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_38c57749[3]));
  AL_DFF_X al_7dcd668a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9868190b[4]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_38c57749[4]));
  AL_DFF_X al_abd0a17c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9868190b[5]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_38c57749[5]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_6a903223 (
    .a(1'b0),
    .o({al_1c02a3cb,open_n2}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6be092bd (
    .a(al_ac3dcbf8[0]),
    .b(1'b1),
    .c(al_1c02a3cb),
    .o({al_ae0d49cd,al_dd86ad38[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3c69ec5 (
    .a(al_ac3dcbf8[1]),
    .b(1'b0),
    .c(al_ae0d49cd),
    .o({al_9df86c79,al_dd86ad38[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_dd382819 (
    .a(al_ac3dcbf8[2]),
    .b(1'b0),
    .c(al_9df86c79),
    .o({al_4f080ff4,al_dd86ad38[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_69231e29 (
    .a(al_ac3dcbf8[3]),
    .b(1'b0),
    .c(al_4f080ff4),
    .o({al_f12d2a54,al_dd86ad38[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_64ebc87c (
    .a(al_ac3dcbf8[4]),
    .b(1'b0),
    .c(al_f12d2a54),
    .o({al_951148c8,al_dd86ad38[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d0dc1a6b (
    .a(al_ac3dcbf8[5]),
    .b(1'b0),
    .c(al_951148c8),
    .o({al_3e63fd9,al_dd86ad38[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d89fb06b (
    .a(al_ac3dcbf8[6]),
    .b(1'b0),
    .c(al_3e63fd9),
    .o({al_19dda09f,al_dd86ad38[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e537e50 (
    .a(al_ac3dcbf8[7]),
    .b(1'b0),
    .c(al_19dda09f),
    .o({al_46b6d0af,al_dd86ad38[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5d65c61d (
    .a(al_ac3dcbf8[8]),
    .b(1'b0),
    .c(al_46b6d0af),
    .o({al_20d13f12,al_dd86ad38[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4431a079 (
    .a(al_ac3dcbf8[9]),
    .b(1'b0),
    .c(al_20d13f12),
    .o({al_3290811f,al_dd86ad38[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7c3f6a55 (
    .a(al_ac3dcbf8[10]),
    .b(1'b0),
    .c(al_3290811f),
    .o({al_e25e65e3,al_dd86ad38[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4ad16480 (
    .a(al_ac3dcbf8[11]),
    .b(1'b0),
    .c(al_e25e65e3),
    .o({al_607f31be,al_dd86ad38[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_86c932ab (
    .a(al_ac3dcbf8[12]),
    .b(1'b0),
    .c(al_607f31be),
    .o({al_b5a71093,al_dd86ad38[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7372f11b (
    .a(al_ac3dcbf8[13]),
    .b(1'b0),
    .c(al_b5a71093),
    .o({al_336a5970,al_dd86ad38[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1a1edd09 (
    .a(al_ac3dcbf8[14]),
    .b(1'b0),
    .c(al_336a5970),
    .o({al_700f8a99,al_dd86ad38[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d84e2848 (
    .a(al_ac3dcbf8[15]),
    .b(1'b0),
    .c(al_700f8a99),
    .o({open_n3,al_dd86ad38[15]}));
  AL_DFF_0 al_52b01358 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_59f1a9e9),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_de12b3ef));
  AL_DFF_0 al_67e559ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_de12b3ef),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_dd6bc6a));
  AL_DFF_X al_69856307 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f6643499),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(tx_retransmit));
  AL_DFF_X al_91dacff9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_stop),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_6b48ce98));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(~A*~(D*C*~B)))"),
    .INIT(32'h0000baaa))
    al_e5874871 (
    .a(tx_status_vector[3]),
    .b(al_1dee2dce[0]),
    .c(al_1dee2dce[1]),
    .d(al_1dee2dce[4]),
    .e(tx_status_vld),
    .o(al_dad1457e));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_27c6d6b6 (
    .a(al_c88c8301),
    .b(al_68462158),
    .o(al_2e1a2363));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_fef0207 (
    .a(al_a09e8e00),
    .b(al_b3be0d17),
    .o(al_3fd53f68));
  AL_DFF_X al_7733ac1c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_data[0]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_251fb86c[0]));
  AL_DFF_X al_27b14679 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_data[1]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_251fb86c[1]));
  AL_DFF_X al_9aa8fe55 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_data[2]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_251fb86c[2]));
  AL_DFF_X al_3d2737bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_data[3]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_251fb86c[3]));
  AL_DFF_X al_d264eb83 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_data[4]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_251fb86c[4]));
  AL_DFF_X al_3b929979 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_data[5]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_251fb86c[5]));
  AL_DFF_X al_49a57d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_data[6]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_251fb86c[6]));
  AL_DFF_X al_46077bc7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_data[7]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_251fb86c[7]));
  AL_DFF_X al_96ff942b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5160c8c2[0]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_data[0]));
  AL_DFF_X al_d2adfb5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5160c8c2[1]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_data[1]));
  AL_DFF_X al_1edc9e1c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5160c8c2[2]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_data[2]));
  AL_DFF_X al_ceb2b8c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5160c8c2[3]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_data[3]));
  AL_DFF_X al_b90d537c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5160c8c2[4]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_data[4]));
  AL_DFF_X al_5bd88b93 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5160c8c2[5]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_data[5]));
  AL_DFF_X al_98ce7d2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5160c8c2[6]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_data[6]));
  AL_DFF_X al_fb89143b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5160c8c2[7]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_data[7]));
  AL_DFF_0 al_3194821d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_a0f12bef[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29842798));
  AL_DFF_0 al_d4d7fd97 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_29842798),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68462158));
  AL_DFF_0 al_b51c20dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_7808e039[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_87773c5e));
  AL_DFF_0 al_108a4db (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_87773c5e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c88c8301));
  AL_DFF_0 al_3008dec (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9b4eaefc[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd1b7e74));
  AL_DFF_0 al_11515b60 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cd1b7e74),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b3be0d17));
  AL_DFF_0 al_5b08f5ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_7808e039[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3cd9a398));
  AL_DFF_0 al_33044622 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_3cd9a398),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a09e8e00));
  AL_DFF_X al_a40fb742 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e2923d0b),
    .en(1'b1),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_4df60ad5));
  AL_DFF_X al_8173e3e1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_2ef0a421),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_88f7ad44));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    al_24d3162f (
    .a(al_ecbdcaf1[0]),
    .b(al_ecbdcaf1[1]),
    .c(al_ecbdcaf1[2]),
    .d(al_ecbdcaf1[3]),
    .o(al_5607a442));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*~C*B*A)"),
    .INIT(32'h00000800))
    al_4691666d (
    .a(al_5607a442),
    .b(al_2e624116[0]),
    .c(al_2e624116[1]),
    .d(al_2e624116[2]),
    .e(al_2e624116[3]),
    .o(al_482a08f7));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_47a27513 (
    .a(al_482a08f7),
    .b(al_d407324e),
    .o(al_8e2f2cc5));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_204d708d (
    .a(al_8e2f2cc5),
    .b(al_ff9a7266),
    .c(al_88f7ad44),
    .o(al_2ef0a421));
  AL_DFF_X al_7965f091 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_379b9322),
    .en(1'b1),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_aa509190));
  AL_DFF_X al_11c9a48c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_aa509190),
    .en(1'b1),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_f766fdfa));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_f32a42c9 (
    .a(al_40258be6),
    .b(al_604d05a2),
    .c(al_76e54a1a),
    .o(al_379b9322));
  AL_DFF_X al_7260aef1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(gmii_rx_vld),
    .en(1'b1),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_49c3c8c7));
  AL_DFF_X al_3bade7b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_49c3c8c7),
    .en(1'b1),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_40258be6));
  AL_DFF_X al_402d11fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f50bd9c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fc6a7e7a));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*~A)"),
    .INIT(16'h0040))
    al_f65a93c6 (
    .a(al_49c3c8c7),
    .b(al_40258be6),
    .c(al_b79f6a7b[0]),
    .d(al_25215c55[1]),
    .o(al_e2923d0b));
  AL_MAP_LUT4 #(
    .EQN("(C*~B*~(~D*A))"),
    .INIT(16'h3010))
    al_1afd96e0 (
    .a(al_e2923d0b),
    .b(al_ff9a7266),
    .c(al_40258be6),
    .d(al_604d05a2),
    .o(al_f50bd9c));
  AL_DFF_X al_cd1ed96a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(gmii_rx_er),
    .en(1'b1),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_755e05f8));
  AL_DFF_X al_74dd52e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_755e05f8),
    .en(1'b1),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_604d05a2));
  AL_DFF_X al_a19e5da5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_604d05a2),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_53de47ce));
  AL_DFF_X al_296046ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_53de47ce),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fc5f2d2a));
  AL_DFF_X al_ce1c44e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_8e2f2cc5),
    .en(1'b1),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_afc1b64));
  AL_DFF_X al_81a4b840 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_afc1b64),
    .en(1'b1),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_76e54a1a));
  AL_DFF_X al_442a695f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b3908a65),
    .en(1'b1),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_d407324e));
  AL_MAP_LUT6 #(
    .EQN("~(~(~D*B)*~(F*~(~E*~C*A)))"),
    .INIT(64'hfffff5fd00cc00cc))
    al_ac9ccaca (
    .a(al_482a08f7),
    .b(al_49c3c8c7),
    .c(al_755e05f8),
    .d(al_40258be6),
    .e(al_604d05a2),
    .f(al_d407324e),
    .o(al_b3908a65));
  AL_DFF_X al_90efb6ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ecbdcaf1[0]),
    .en(1'b1),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_2e624116[0]));
  AL_DFF_X al_1dfb8f94 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ecbdcaf1[1]),
    .en(1'b1),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_2e624116[1]));
  AL_DFF_X al_977a9e43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ecbdcaf1[2]),
    .en(1'b1),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_2e624116[2]));
  AL_DFF_X al_8c38fc42 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ecbdcaf1[3]),
    .en(1'b1),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_2e624116[3]));
  AL_DFF_X al_c41a1e51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_2e624116[0]),
    .en(1'b1),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_d286f1cd[0]));
  AL_DFF_X al_b6d5b3f3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_2e624116[1]),
    .en(1'b1),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_d286f1cd[1]));
  AL_DFF_X al_22cf5b7c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_2e624116[2]),
    .en(1'b1),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_d286f1cd[2]));
  AL_DFF_X al_5492b5e1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_2e624116[3]),
    .en(1'b1),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_d286f1cd[3]));
  AL_DFF_X al_b890aec3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_d286f1cd[0]),
    .en(1'b1),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_62f364a9[0]));
  AL_DFF_X al_1a6b1341 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_d286f1cd[1]),
    .en(1'b1),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_62f364a9[1]));
  AL_DFF_X al_d30cd802 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_d286f1cd[2]),
    .en(1'b1),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_62f364a9[2]));
  AL_DFF_X al_85b9f768 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_d286f1cd[3]),
    .en(1'b1),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_62f364a9[3]));
  AL_DFF_X al_358a0deb (
    .ar(al_d407324e),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_d9ec2230),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b79f6a7b[0]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_fd4834d9 (
    .a(al_40258be6),
    .b(al_b79f6a7b[0]),
    .o(al_d9ec2230));
  AL_DFF_X al_f9a17bc9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(gmii_rxd[0]),
    .en(1'b1),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_ecbdcaf1[0]));
  AL_DFF_X al_319f3fd9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(gmii_rxd[1]),
    .en(1'b1),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_ecbdcaf1[1]));
  AL_DFF_X al_9c013c6b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(gmii_rxd[2]),
    .en(1'b1),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_ecbdcaf1[2]));
  AL_DFF_X al_483e69ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(gmii_rxd[3]),
    .en(1'b1),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_ecbdcaf1[3]));
  AL_DFF_X al_d76ed390 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(gmii_rxd[4]),
    .en(1'b1),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_ecbdcaf1[4]));
  AL_DFF_X al_6b6ec17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(gmii_rxd[5]),
    .en(1'b1),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_ecbdcaf1[5]));
  AL_DFF_X al_1a4e9b67 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(gmii_rxd[6]),
    .en(1'b1),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_ecbdcaf1[6]));
  AL_DFF_X al_e98dc4d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(gmii_rxd[7]),
    .en(1'b1),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_ecbdcaf1[7]));
  AL_DFF_X al_5855ed95 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(gmii_col),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_7c904594));
  AL_DFF_X al_a13f5ebe (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_7c904594),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_f785157a));
  AL_DFF_X al_7c53e4e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d75651de),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_b4b52182));
  AL_DFF_X al_cf81f2fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b4b52182),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_44e126e5));
  AL_DFF_X al_554617ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_52e770ef),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_3dc7e6d6));
  AL_DFF_X al_1bfc3162 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_25291b5c),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_1a7bad30));
  AL_DFF_X al_77444f13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1cbba6e6),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_e5091a32));
  AL_DFF_X al_1e3b5ca8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_372f5c11),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_5d53f279));
  AL_DFF_X al_10fe28ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_8aa33695),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_26f70e9a));
  AL_DFF_X al_873bb722 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_26f70e9a),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_186c00a8));
  AL_DFF_X al_d4a708bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1f250659),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_3c343df4));
  AL_DFF_X al_ec181f13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_3c343df4),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_21c59f1));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*~(D)*~(E)+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*D*~(E)+~((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))*D*E+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*D*E)"),
    .INIT(32'hff00caca))
    al_28f1a767 (
    .a(al_78b1b46e[0]),
    .b(al_78b1b46e[4]),
    .c(al_5d53f279),
    .d(al_b25edb3[0]),
    .e(al_25215c55[1]),
    .o(al_fbc4ef28[0]));
  AL_MAP_LUT5 #(
    .EQN("~(~C*~(D*~B)*~(~E*A))"),
    .INIT(32'hf3f0fbfa))
    al_e433677a (
    .a(al_22c188eb),
    .b(al_a6f148e9),
    .c(al_4a547188),
    .d(al_fbc4ef28[0]),
    .e(al_a49d6a86),
    .o(al_5bef7ee6[0]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*~(D)*~(E)+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*D*~(E)+~((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))*D*E+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*D*E)"),
    .INIT(32'hff00caca))
    al_efaa3061 (
    .a(al_78b1b46e[1]),
    .b(al_78b1b46e[5]),
    .c(al_5d53f279),
    .d(al_b25edb3[1]),
    .e(al_25215c55[1]),
    .o(al_fbc4ef28[1]));
  AL_MAP_LUT5 #(
    .EQN("~(~C*~(D*~B)*~(~E*A))"),
    .INIT(32'hf3f0fbfa))
    al_8b992d91 (
    .a(al_22c188eb),
    .b(al_a6f148e9),
    .c(al_4a547188),
    .d(al_fbc4ef28[1]),
    .e(al_a49d6a86),
    .o(al_5bef7ee6[1]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*~(D)*~(E)+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*D*~(E)+~((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))*D*E+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*D*E)"),
    .INIT(32'hff00caca))
    al_6f238a7c (
    .a(al_78b1b46e[2]),
    .b(al_78b1b46e[6]),
    .c(al_5d53f279),
    .d(al_b25edb3[2]),
    .e(al_25215c55[1]),
    .o(al_fbc4ef28[2]));
  AL_MAP_LUT5 #(
    .EQN("~(~C*~(D*~B)*~(~E*A))"),
    .INIT(32'hf3f0fbfa))
    al_a01fe4a3 (
    .a(al_22c188eb),
    .b(al_a6f148e9),
    .c(al_4a547188),
    .d(al_fbc4ef28[2]),
    .e(al_a49d6a86),
    .o(al_5bef7ee6[2]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*~(D)*~(E)+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*D*~(E)+~((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))*D*E+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*D*E)"),
    .INIT(32'hff00caca))
    al_bab52160 (
    .a(al_78b1b46e[3]),
    .b(al_78b1b46e[7]),
    .c(al_5d53f279),
    .d(al_b25edb3[3]),
    .e(al_25215c55[1]),
    .o(al_fbc4ef28[3]));
  AL_MAP_LUT5 #(
    .EQN("~(~C*~(D*~B)*~(~E*A))"),
    .INIT(32'hf3f0fbfa))
    al_de1f00ea (
    .a(al_22c188eb),
    .b(al_a6f148e9),
    .c(al_4a547188),
    .d(al_fbc4ef28[3]),
    .e(al_a49d6a86),
    .o(al_5bef7ee6[3]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_3aa22c2c (
    .a(al_20d4193c[0]),
    .b(al_20d4193c[1]),
    .c(al_20d4193c[2]),
    .o(al_9b6b0ae2));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    al_4bb06bfe (
    .a(al_26f70e9a),
    .b(al_186c00a8),
    .c(al_3dc7e6d6),
    .d(al_25215c55[1]),
    .o(al_72ac780f));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    al_a8d8a9ca (
    .a(al_72ac780f),
    .b(al_96252128[0]),
    .c(al_96252128[1]),
    .d(al_96252128[2]),
    .e(al_96252128[3]),
    .o(al_7978050f));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    al_b1bfb4fc (
    .a(al_7978050f),
    .b(al_9b6b0ae2),
    .c(al_20d4193c[3]),
    .o(al_22c188eb));
  AL_MAP_LUT6 #(
    .EQN("(~A*~((~E*~D)*~((~C*~B))*~(F)+(~E*~D)*(~C*~B)*~(F)+~((~E*~D))*(~C*~B)*F+(~E*~D)*(~C*~B)*F))"),
    .INIT(64'h5454545455555500))
    al_43a4a413 (
    .a(al_bb1dc6ea),
    .b(al_d2863baf[3]),
    .c(al_d2863baf[5]),
    .d(al_d2863baf[7]),
    .e(al_d2863baf[11]),
    .f(al_25215c55[1]),
    .o(al_a6f148e9));
  AL_MAP_LUT6 #(
    .EQN("~(~C*~(F*E*~B)*~(~D*A))"),
    .INIT(64'hf3fbf0faf0faf0fa))
    al_fe5c1a08 (
    .a(al_22c188eb),
    .b(al_a6f148e9),
    .c(al_4a547188),
    .d(al_a49d6a86),
    .e(al_b25edb3[4]),
    .f(al_25215c55[1]),
    .o(al_5bef7ee6[4]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_44acd4b (
    .a(al_a59c7c46[0]),
    .b(al_a59c7c46[1]),
    .c(al_a59c7c46[2]),
    .d(al_a59c7c46[3]),
    .o(al_f8bfe558));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*A)"),
    .INIT(8'hf7))
    al_ec2a07c7 (
    .a(al_f8bfe558),
    .b(al_9b6b0ae2),
    .c(al_20d4193c[3]),
    .o(al_bb1dc6ea));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_7c0b1a10 (
    .a(al_b4b52182),
    .b(al_44e126e5),
    .c(al_25215c55[1]),
    .o(al_a49d6a86));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_9ad77cbd (
    .a(al_f8bfe558),
    .b(al_a49d6a86),
    .o(al_4a547188));
  AL_MAP_LUT6 #(
    .EQN("~(~(F*E*~C*~B)*~(~D*A))"),
    .INIT(64'h03ab00aa00aa00aa))
    al_39527f97 (
    .a(al_22c188eb),
    .b(al_a6f148e9),
    .c(al_4a547188),
    .d(al_a49d6a86),
    .e(al_b25edb3[5]),
    .f(al_25215c55[1]),
    .o(al_5bef7ee6[5]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F*E*~C*~B)*~(~D*A))"),
    .INIT(64'h03ab00aa00aa00aa))
    al_107766cc (
    .a(al_22c188eb),
    .b(al_a6f148e9),
    .c(al_4a547188),
    .d(al_a49d6a86),
    .e(al_b25edb3[6]),
    .f(al_25215c55[1]),
    .o(al_5bef7ee6[6]));
  AL_MAP_LUT6 #(
    .EQN("~(~(F*E*~C*~B)*~(~D*A))"),
    .INIT(64'h03ab00aa00aa00aa))
    al_13e91700 (
    .a(al_22c188eb),
    .b(al_a6f148e9),
    .c(al_4a547188),
    .d(al_a49d6a86),
    .e(al_b25edb3[7]),
    .f(al_25215c55[1]),
    .o(al_5bef7ee6[7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_22af5dd7 (
    .a(al_26f70e9a),
    .b(al_186c00a8),
    .c(al_25215c55[1]),
    .o(al_52e770ef));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(D*~B*~(~E*~C)))"),
    .INIT(32'hbbaabaaa))
    al_54f4083b (
    .a(al_22c188eb),
    .b(al_a6f148e9),
    .c(al_f8bfe558),
    .d(al_52e770ef),
    .e(al_d75651de),
    .o(al_25291b5c));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_b0036451 (
    .a(al_3c343df4),
    .b(al_21c59f1),
    .c(al_25215c55[1]),
    .o(al_cd3fff34));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(~(~E*~C)*~(D*~B)))"),
    .INIT(32'h11001505))
    al_60921a02 (
    .a(al_22c188eb),
    .b(al_a6f148e9),
    .c(al_f8bfe558),
    .d(al_cd3fff34),
    .e(al_d75651de),
    .o(al_1cbba6e6));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*A))"),
    .INIT(8'h0d))
    al_3ceaa7a0 (
    .a(al_26f70e9a),
    .b(al_186c00a8),
    .c(al_5d53f279),
    .o(al_372f5c11));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    al_88d1b0e4 (
    .a(al_7978050f),
    .b(al_72ac780f),
    .c(al_96252128[0]),
    .o(al_dc435ff2[0]));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~B*(D@C)))"),
    .INIT(16'h5445))
    al_912dc6ce (
    .a(al_7978050f),
    .b(al_72ac780f),
    .c(al_96252128[0]),
    .d(al_96252128[1]),
    .o(al_dc435ff2[1]));
  AL_MAP_LUT5 #(
    .EQN("~(~A*(~((~C*~B))*~(D)*~(E)+(~C*~B)*~(D)*~(E)+(~C*~B)*D*~(E)+~((~C*~B))*~(D)*E+(~C*~B)*D*E))"),
    .INIT(32'hfeabfeaa))
    al_b6517887 (
    .a(al_72ac780f),
    .b(al_96252128[0]),
    .c(al_96252128[1]),
    .d(al_96252128[2]),
    .e(al_96252128[3]),
    .o(al_dc435ff2[2]));
  AL_MAP_LUT6 #(
    .EQN("~(~(E*~(~D*~C*~B))*~(F)*~(A)+~(E*~(~D*~C*~B))*F*~(A)+~(~(E*~(~D*~C*~B)))*F*A+~(E*~(~D*~C*~B))*F*A)"),
    .INIT(64'h55540000fffeaaaa))
    al_284e583b (
    .a(al_72ac780f),
    .b(al_96252128[0]),
    .c(al_96252128[1]),
    .d(al_96252128[2]),
    .e(al_96252128[3]),
    .f(al_25215c55[1]),
    .o(al_dc435ff2[3]));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_3a06eded (
    .a(al_22c188eb),
    .b(al_25dd3b31),
    .c(al_20d4193c[0]),
    .o(al_ee96b553[0]));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(~C*A)))"),
    .INIT(16'h3102))
    al_e7581737 (
    .a(al_22c188eb),
    .b(al_25dd3b31),
    .c(al_20d4193c[0]),
    .d(al_20d4193c[1]),
    .o(al_ee96b553[1]));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    al_77b4c07e (
    .a(al_52e770ef),
    .b(al_7c904594),
    .c(al_f785157a),
    .d(al_9b4eaefc[2]),
    .o(al_25dd3b31));
  AL_MAP_LUT6 #(
    .EQN("((E@(~D*~C*A))*~(F)*~(B)+(E@(~D*~C*A))*F*~(B)+~((E@(~D*~C*A)))*F*B+(E@(~D*~C*A))*F*B)"),
    .INIT(64'hfffdccce33310002))
    al_92d48600 (
    .a(al_22c188eb),
    .b(al_25dd3b31),
    .c(al_20d4193c[0]),
    .d(al_20d4193c[1]),
    .e(al_20d4193c[2]),
    .f(al_25215c55[1]),
    .o(al_ee96b553[2]));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*~(C*A))*~(E)*~(B)+~(D*~(C*A))*E*~(B)+~(~(D*~(C*A)))*E*B+~(D*~(C*A))*E*B)"),
    .INIT(32'h1300dfcc))
    al_d9650e39 (
    .a(al_7978050f),
    .b(al_25dd3b31),
    .c(al_9b6b0ae2),
    .d(al_20d4193c[3]),
    .e(al_25215c55[1]),
    .o(al_ee96b553[3]));
  AL_MAP_LUT3 #(
    .EQN("(~A*(C@B))"),
    .INIT(8'h14))
    al_e4770a55 (
    .a(al_8edce7a2),
    .b(al_4a547188),
    .c(al_a59c7c46[0]),
    .o(al_95650af7[0]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D@(~C*B)))"),
    .INIT(16'h5104))
    al_82726a84 (
    .a(al_8edce7a2),
    .b(al_4a547188),
    .c(al_a59c7c46[0]),
    .d(al_a59c7c46[1]),
    .o(al_95650af7[1]));
  AL_MAP_LUT6 #(
    .EQN("(F*~E*D*C*B*~A)"),
    .INIT(64'h0000400000000000))
    al_d504f3a6 (
    .a(al_52e770ef),
    .b(al_cd3fff34),
    .c(al_a49d6a86),
    .d(al_7c904594),
    .e(al_f785157a),
    .f(al_9b4eaefc[2]),
    .o(al_8edce7a2));
  AL_MAP_LUT6 #(
    .EQN("((E@(~D*~C*B))*~(F)*~(A)+(E@(~D*~C*B))*F*~(A)+~((E@(~D*~C*B)))*F*A+(E@(~D*~C*B))*F*A)"),
    .INIT(64'hfffbaaae55510004))
    al_52657787 (
    .a(al_8edce7a2),
    .b(al_4a547188),
    .c(al_a59c7c46[0]),
    .d(al_a59c7c46[1]),
    .e(al_a59c7c46[2]),
    .f(al_25215c55[1]),
    .o(al_95650af7[2]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_c1f5166f (
    .a(al_a59c7c46[0]),
    .b(al_a59c7c46[1]),
    .c(al_a59c7c46[2]),
    .o(al_674bc53d));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*~(~C*B))*~(E)*~(A)+~(D*~(~C*B))*E*~(A)+~(~(D*~(~C*B)))*E*A+~(D*~(~C*B))*E*A)"),
    .INIT(32'h5100fbaa))
    al_813132be (
    .a(al_8edce7a2),
    .b(al_674bc53d),
    .c(al_a49d6a86),
    .d(al_a59c7c46[3]),
    .e(al_25215c55[1]),
    .o(al_95650af7[3]));
  AL_DFF_X al_1056349b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b25edb3[0]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_78b1b46e[0]));
  AL_DFF_X al_8aa94dc9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b25edb3[1]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_78b1b46e[1]));
  AL_DFF_X al_6b1b5d89 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b25edb3[2]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_78b1b46e[2]));
  AL_DFF_X al_1d3b7465 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b25edb3[3]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_78b1b46e[3]));
  AL_DFF_X al_5fe2036d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b25edb3[4]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_78b1b46e[4]));
  AL_DFF_X al_67a5c223 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b25edb3[5]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_78b1b46e[5]));
  AL_DFF_X al_7ec057e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b25edb3[6]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_78b1b46e[6]));
  AL_DFF_X al_21aa1aba (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b25edb3[7]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_78b1b46e[7]));
  AL_DFF_X al_60a4cb67 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5bef7ee6[0]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_bb772f98[0]));
  AL_DFF_X al_55183cde (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5bef7ee6[1]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_bb772f98[1]));
  AL_DFF_X al_c235bb63 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5bef7ee6[2]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_bb772f98[2]));
  AL_DFF_X al_5a211588 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5bef7ee6[3]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_bb772f98[3]));
  AL_DFF_X al_26b6b40e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5bef7ee6[4]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_bb772f98[4]));
  AL_DFF_X al_fe533efe (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5bef7ee6[5]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_bb772f98[5]));
  AL_DFF_X al_74305ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5bef7ee6[6]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_bb772f98[6]));
  AL_DFF_X al_fa4512c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5bef7ee6[7]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_bb772f98[7]));
  AL_DFF_X al_622545d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_dc435ff2[0]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_96252128[0]));
  AL_DFF_X al_ad6f62a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_dc435ff2[1]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_96252128[1]));
  AL_DFF_X al_6e6cc291 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_dc435ff2[2]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_96252128[2]));
  AL_DFF_X al_65a4d32f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_dc435ff2[3]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_96252128[3]));
  AL_DFF_X al_bf5f6743 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ee96b553[0]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_20d4193c[0]));
  AL_DFF_X al_5ddd78e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ee96b553[1]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_20d4193c[1]));
  AL_DFF_X al_e2dc3752 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ee96b553[2]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_20d4193c[2]));
  AL_DFF_X al_e6fd2871 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ee96b553[3]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_20d4193c[3]));
  AL_DFF_X al_bac0c66 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_95650af7[0]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_a59c7c46[0]));
  AL_DFF_X al_c4e1e590 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_95650af7[1]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_a59c7c46[1]));
  AL_DFF_X al_83b314d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_95650af7[2]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_a59c7c46[2]));
  AL_DFF_X al_db751ffa (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_95650af7[3]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_a59c7c46[3]));
  AL_DFF_X al_a666aba9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_bb1dc6ea),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_d2863baf[0]));
  AL_DFF_X al_dbd22c6c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d2863baf[8]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_d2863baf[9]));
  AL_DFF_X al_3963f8ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d2863baf[9]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_d2863baf[10]));
  AL_DFF_X al_37e2565f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d2863baf[10]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_d2863baf[11]));
  AL_DFF_X al_89cbc351 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d2863baf[0]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_d2863baf[1]));
  AL_DFF_X al_b6db5f5a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d2863baf[1]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_d2863baf[2]));
  AL_DFF_X al_966b3545 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d2863baf[2]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_d2863baf[3]));
  AL_DFF_X al_f9098a67 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d2863baf[3]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_d2863baf[4]));
  AL_DFF_X al_eff0f77 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d2863baf[4]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_d2863baf[5]));
  AL_DFF_X al_37dc87df (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d2863baf[5]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_d2863baf[6]));
  AL_DFF_X al_76cc92d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d2863baf[6]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_d2863baf[7]));
  AL_DFF_X al_40272ffa (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d2863baf[7]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_d2863baf[8]));
  AL_DFF_X al_656abf38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_96e5a141[0]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_b25edb3[0]));
  AL_DFF_X al_7f886ac7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_96e5a141[1]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_b25edb3[1]));
  AL_DFF_X al_ddfca1e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_96e5a141[2]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_b25edb3[2]));
  AL_DFF_X al_f46abc38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_96e5a141[3]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_b25edb3[3]));
  AL_DFF_X al_dd5e636a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_96e5a141[4]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_b25edb3[4]));
  AL_DFF_X al_33ac9d66 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_96e5a141[5]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_b25edb3[5]));
  AL_DFF_X al_2eb5c816 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_96e5a141[6]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_b25edb3[6]));
  AL_DFF_X al_4f8a7c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_96e5a141[7]),
    .en(gmii_tx_clken),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_b25edb3[7]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*~(D)*~(E)+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*D*~(E)+~((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))*D*E+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*D*E)"),
    .INIT(32'hff00caca))
    al_19cd6d50 (
    .a(al_d286f1cd[0]),
    .b(al_62f364a9[0]),
    .c(al_88f7ad44),
    .d(al_ecbdcaf1[0]),
    .e(al_25215c55[1]),
    .o(al_fa90a029[0]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*~(D)*~(E)+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*D*~(E)+~((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))*D*E+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*D*E)"),
    .INIT(32'hff00caca))
    al_9fcda57e (
    .a(al_d286f1cd[1]),
    .b(al_62f364a9[1]),
    .c(al_88f7ad44),
    .d(al_ecbdcaf1[1]),
    .e(al_25215c55[1]),
    .o(al_fa90a029[1]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*~(D)*~(E)+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*D*~(E)+~((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))*D*E+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*D*E)"),
    .INIT(32'hff00caca))
    al_9d68b565 (
    .a(al_d286f1cd[2]),
    .b(al_62f364a9[2]),
    .c(al_88f7ad44),
    .d(al_ecbdcaf1[2]),
    .e(al_25215c55[1]),
    .o(al_fa90a029[2]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*~(D)*~(E)+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*D*~(E)+~((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))*D*E+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*D*E)"),
    .INIT(32'hff00caca))
    al_f2e93ad4 (
    .a(al_d286f1cd[3]),
    .b(al_62f364a9[3]),
    .c(al_88f7ad44),
    .d(al_ecbdcaf1[3]),
    .e(al_25215c55[1]),
    .o(al_fa90a029[3]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*~(D)*~(E)+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*D*~(E)+~((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))*D*E+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*D*E)"),
    .INIT(32'hff00caca))
    al_8965386 (
    .a(al_2e624116[0]),
    .b(al_d286f1cd[0]),
    .c(al_88f7ad44),
    .d(al_ecbdcaf1[4]),
    .e(al_25215c55[1]),
    .o(al_fa90a029[4]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*~(D)*~(E)+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*D*~(E)+~((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))*D*E+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*D*E)"),
    .INIT(32'hff00caca))
    al_96f390e2 (
    .a(al_2e624116[1]),
    .b(al_d286f1cd[1]),
    .c(al_88f7ad44),
    .d(al_ecbdcaf1[5]),
    .e(al_25215c55[1]),
    .o(al_fa90a029[5]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*~(D)*~(E)+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*D*~(E)+~((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))*D*E+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*D*E)"),
    .INIT(32'hff00caca))
    al_9d9eec73 (
    .a(al_2e624116[2]),
    .b(al_d286f1cd[2]),
    .c(al_88f7ad44),
    .d(al_ecbdcaf1[6]),
    .e(al_25215c55[1]),
    .o(al_fa90a029[6]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*~(D)*~(E)+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*D*~(E)+~((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))*D*E+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*D*E)"),
    .INIT(32'hff00caca))
    al_1ba72617 (
    .a(al_2e624116[3]),
    .b(al_d286f1cd[3]),
    .c(al_88f7ad44),
    .d(al_ecbdcaf1[7]),
    .e(al_25215c55[1]),
    .o(al_fa90a029[7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    al_26ecc3bd (
    .a(al_49c3c8c7),
    .b(al_fc6a7e7a),
    .c(al_25215c55[1]),
    .o(al_46f5ce71));
  AL_MAP_LUT4 #(
    .EQN("(~D*~A*~(C*B))"),
    .INIT(16'h0015))
    al_739e5a69 (
    .a(al_53de47ce),
    .b(al_fc5f2d2a),
    .c(al_88f7ad44),
    .d(al_f766fdfa),
    .o(al_ed888342));
  AL_MAP_LUT6 #(
    .EQN("(~(A*~(~E*D*C))*~(B)*~(F)+~(A*~(~E*D*C))*B*~(F)+~(~(A*~(~E*D*C)))*B*F+~(A*~(~E*D*C))*B*F)"),
    .INIT(64'hcccccccc5555f555))
    al_30ba6faf (
    .a(al_ed888342),
    .b(al_755e05f8),
    .c(al_40258be6),
    .d(al_604d05a2),
    .e(al_76e54a1a),
    .f(al_25215c55[1]),
    .o(al_89fbca82));
  AL_DFF_X al_818403ad (
    .ar(1'b0),
    .as(reset),
    .clk(s_axi_aclk),
    .d(1'b0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59850dc4));
  AL_DFF_X al_763dd809 (
    .ar(1'b0),
    .as(reset),
    .clk(s_axi_aclk),
    .d(al_59850dc4),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_90484227));
  AL_DFF_X al_a9d62e8f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_90484227),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f17b93eb));
  AL_DFF_X al_a559606c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_f517c689),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_81344cef));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_d68c8db6 (
    .a(al_90484227),
    .b(al_f17b93eb),
    .o(al_f517c689));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_50bb8698 (
    .a(reset),
    .b(al_a0f12bef[0]),
    .o(al_1e2edecf));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_cf5c85b2 (
    .a(al_251fb86c[0]),
    .b(al_b984f6c1),
    .c(al_45ed4524[0]),
    .o(al_5db4ba74[0]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_7a1829c1 (
    .a(al_251fb86c[1]),
    .b(al_b984f6c1),
    .c(al_45ed4524[1]),
    .o(al_5db4ba74[1]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_d2fb3e5a (
    .a(al_251fb86c[2]),
    .b(al_b984f6c1),
    .c(al_45ed4524[2]),
    .o(al_5db4ba74[2]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_577fa023 (
    .a(al_251fb86c[3]),
    .b(al_b984f6c1),
    .c(al_45ed4524[3]),
    .o(al_5db4ba74[3]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_aa4564c8 (
    .a(al_251fb86c[4]),
    .b(al_b984f6c1),
    .c(al_45ed4524[4]),
    .o(al_5db4ba74[4]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_75ce4c89 (
    .a(al_251fb86c[5]),
    .b(al_b984f6c1),
    .c(al_45ed4524[5]),
    .o(al_5db4ba74[5]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_2ff29525 (
    .a(al_251fb86c[6]),
    .b(al_b984f6c1),
    .c(al_45ed4524[6]),
    .o(al_5db4ba74[6]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_f5044922 (
    .a(al_251fb86c[7]),
    .b(al_b984f6c1),
    .c(al_45ed4524[7]),
    .o(al_5db4ba74[7]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_720676a4 (
    .a(reset),
    .b(al_9b4eaefc[0]),
    .o(al_6d2cc211));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_a85e2f36 (
    .a(al_b984f6c1),
    .b(al_9b4eaefc[3]),
    .o(al_aa427d37));
  AL_DFF_X al_336c1a01 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_1b903e6a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6b181c0));
  AL_MAP_LUT6 #(
    .EQN("(B*A*~(F@D)*~(E@C))"),
    .INIT(64'h8000080000800008))
    al_f74ff5ba (
    .a(al_35f01e82),
    .b(al_fd6c10a8),
    .c(al_ddeffb0f[4]),
    .d(al_ddeffb0f[5]),
    .e(al_4096d0c7[4]),
    .f(al_4096d0c7[5]),
    .o(al_5bf34257));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*(D@A))"),
    .INIT(16'h0102))
    al_c38877e8 (
    .a(al_5bf34257),
    .b(al_37d9882e),
    .c(al_81344cef),
    .d(al_6b181c0),
    .o(al_1b903e6a));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    al_2a93a5b1 (
    .a(al_ddeffb0f[2]),
    .b(al_ddeffb0f[3]),
    .c(al_4096d0c7[2]),
    .d(al_4096d0c7[3]),
    .o(al_35f01e82));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    al_19daf9b3 (
    .a(al_ddeffb0f[0]),
    .b(al_ddeffb0f[1]),
    .c(al_4096d0c7[0]),
    .d(al_4096d0c7[1]),
    .o(al_fd6c10a8));
  AL_DFF_X al_84b2efca (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_90591ccb),
    .en(1'b1),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_8587a543));
  AL_MAP_LUT5 #(
    .EQN("~(~(~(E*~D)*B)*~(C*A))"),
    .INIT(32'heca0ecec))
    al_c52c23b3 (
    .a(al_fd9c8287),
    .b(al_8587a543),
    .c(al_523025ae[0]),
    .d(al_2b48f483),
    .e(al_841146bf),
    .o(al_90591ccb));
  AL_DFF_X al_a9ba1a3d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_86d0105a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ddeffb0f[0]));
  AL_DFF_X al_cf97ecc (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_1c8c2124),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ddeffb0f[1]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_bdd32cf1 (
    .a(al_5bf34257),
    .b(al_81344cef),
    .o(al_4c800f86));
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'h28))
    al_6631ba0e (
    .a(al_4c800f86),
    .b(al_ddeffb0f[0]),
    .c(al_ddeffb0f[1]),
    .o(al_1c8c2124));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_3eab2abc (
    .a(al_4c800f86),
    .b(al_ddeffb0f[0]),
    .o(al_86d0105a));
  AL_MAP_LUT4 #(
    .EQN("(A*(D@(C*B)))"),
    .INIT(16'h2a80))
    al_65f30970 (
    .a(al_4c800f86),
    .b(al_ddeffb0f[0]),
    .c(al_ddeffb0f[1]),
    .d(al_ddeffb0f[2]),
    .o(al_adafc833));
  AL_MAP_LUT5 #(
    .EQN("(A*(E@(D*C*B)))"),
    .INIT(32'h2aaa8000))
    al_4b6b2dda (
    .a(al_4c800f86),
    .b(al_ddeffb0f[0]),
    .c(al_ddeffb0f[1]),
    .d(al_ddeffb0f[2]),
    .e(al_ddeffb0f[3]),
    .o(al_fb0d0f97));
  AL_DFF_X al_58e76ebb (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_adafc833),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ddeffb0f[2]));
  AL_MAP_LUT6 #(
    .EQN("(A*(F@(E*D*C*B)))"),
    .INIT(64'h2aaaaaaa80000000))
    al_a6ef3d7 (
    .a(al_4c800f86),
    .b(al_ddeffb0f[0]),
    .c(al_ddeffb0f[1]),
    .d(al_ddeffb0f[2]),
    .e(al_ddeffb0f[3]),
    .f(al_ddeffb0f[4]),
    .o(al_7fbfd2c7));
  AL_MAP_LUT6 #(
    .EQN("(F@(E*D*C*B*A))"),
    .INIT(64'h7fffffff80000000))
    al_b8050c0 (
    .a(al_ddeffb0f[0]),
    .b(al_ddeffb0f[1]),
    .c(al_ddeffb0f[2]),
    .d(al_ddeffb0f[3]),
    .e(al_ddeffb0f[4]),
    .f(al_ddeffb0f[5]),
    .o(al_58820abe[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_e53c83e6 (
    .a(al_4c800f86),
    .b(al_58820abe[5]),
    .o(al_63bd33e6));
  AL_DFF_X al_67e0304c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_fb0d0f97),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ddeffb0f[3]));
  AL_DFF_X al_2b8a3861 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_7fbfd2c7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ddeffb0f[4]));
  AL_DFF_X al_5955e9e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_63bd33e6),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ddeffb0f[5]));
  AL_DFF_X al_48b5500e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_a584e1fd),
    .en(1'b1),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(s_axi_arready));
  AL_DFF_X al_7aac7f3f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_bf676c3e),
    .en(1'b1),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(s_axi_bvalid));
  AL_DFF_X al_26390d2e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_1d703c48),
    .en(1'b1),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(s_axi_rvalid));
  AL_DFF_X al_9fc4226 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_dbd330f5),
    .en(1'b1),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(s_axi_wready));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*~B*A)"),
    .INIT(32'h00000020))
    al_3dd4b95 (
    .a(al_cf696ef0),
    .b(al_13660933[4]),
    .c(al_13660933[5]),
    .d(al_13660933[6]),
    .e(al_13660933[7]),
    .o(al_291f5813));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_31a280d3 (
    .a(al_291f5813),
    .b(s_axi_wdata[0]),
    .o(al_624c8b6f));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    al_957254cf (
    .a(al_cf696ef0),
    .b(al_13660933[4]),
    .c(al_13660933[5]),
    .d(al_13660933[6]),
    .e(al_13660933[7]),
    .o(al_c3d9ce92));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_873a9dad (
    .a(al_c3d9ce92),
    .b(s_axi_wdata[0]),
    .o(al_e7647890));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_172ff4ba (
    .a(al_81344cef),
    .b(al_9b4eaefc[0]),
    .o(al_1b655917));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_2f25044c (
    .a(al_ad19785e),
    .b(al_35a8bfef),
    .c(pause_source_addr[0]),
    .d(s_axi_wdata[0]),
    .e(al_868a1cad[0]),
    .o(al_238a702c[0]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_17815f3e (
    .a(al_ad19785e),
    .b(al_35a8bfef),
    .c(pause_source_addr[10]),
    .d(s_axi_wdata[10]),
    .e(al_868a1cad[10]),
    .o(al_238a702c[10]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_6fc023c2 (
    .a(al_ad19785e),
    .b(al_35a8bfef),
    .c(pause_source_addr[11]),
    .d(s_axi_wdata[11]),
    .e(al_868a1cad[11]),
    .o(al_238a702c[11]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_f25df407 (
    .a(al_ad19785e),
    .b(al_35a8bfef),
    .c(pause_source_addr[12]),
    .d(s_axi_wdata[12]),
    .e(al_868a1cad[12]),
    .o(al_238a702c[12]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_889dc374 (
    .a(al_ad19785e),
    .b(al_35a8bfef),
    .c(pause_source_addr[13]),
    .d(s_axi_wdata[13]),
    .e(al_868a1cad[13]),
    .o(al_238a702c[13]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_a77c3ad4 (
    .a(al_ad19785e),
    .b(al_35a8bfef),
    .c(pause_source_addr[14]),
    .d(s_axi_wdata[14]),
    .e(al_868a1cad[14]),
    .o(al_238a702c[14]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_d73efc9 (
    .a(al_ad19785e),
    .b(al_35a8bfef),
    .c(pause_source_addr[15]),
    .d(s_axi_wdata[15]),
    .e(al_868a1cad[15]),
    .o(al_238a702c[15]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_333991d2 (
    .a(al_ad19785e),
    .b(al_35a8bfef),
    .c(pause_source_addr[16]),
    .d(s_axi_wdata[16]),
    .e(al_868a1cad[16]),
    .o(al_238a702c[16]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_43069dbd (
    .a(al_ad19785e),
    .b(al_35a8bfef),
    .c(pause_source_addr[17]),
    .d(s_axi_wdata[17]),
    .e(al_868a1cad[17]),
    .o(al_238a702c[17]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_de486d3c (
    .a(al_ad19785e),
    .b(al_35a8bfef),
    .c(pause_source_addr[18]),
    .d(s_axi_wdata[18]),
    .e(al_868a1cad[18]),
    .o(al_238a702c[18]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_213fdfeb (
    .a(al_ad19785e),
    .b(al_35a8bfef),
    .c(pause_source_addr[19]),
    .d(s_axi_wdata[19]),
    .e(al_868a1cad[19]),
    .o(al_238a702c[19]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_a1993433 (
    .a(al_ad19785e),
    .b(al_35a8bfef),
    .c(pause_source_addr[1]),
    .d(s_axi_wdata[1]),
    .e(al_868a1cad[1]),
    .o(al_238a702c[1]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_e540ae2e (
    .a(al_ad19785e),
    .b(al_35a8bfef),
    .c(pause_source_addr[20]),
    .d(s_axi_wdata[20]),
    .e(al_868a1cad[20]),
    .o(al_238a702c[20]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_f0d88652 (
    .a(al_ad19785e),
    .b(al_35a8bfef),
    .c(pause_source_addr[21]),
    .d(s_axi_wdata[21]),
    .e(al_868a1cad[21]),
    .o(al_238a702c[21]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_65267d2d (
    .a(al_ad19785e),
    .b(al_35a8bfef),
    .c(pause_source_addr[22]),
    .d(s_axi_wdata[22]),
    .e(al_868a1cad[22]),
    .o(al_238a702c[22]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_338f4b85 (
    .a(al_ad19785e),
    .b(al_35a8bfef),
    .c(pause_source_addr[23]),
    .d(s_axi_wdata[23]),
    .e(al_868a1cad[23]),
    .o(al_238a702c[23]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_f773555 (
    .a(al_ad19785e),
    .b(al_35a8bfef),
    .c(pause_source_addr[24]),
    .d(s_axi_wdata[24]),
    .e(al_868a1cad[24]),
    .o(al_238a702c[24]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_b41318dd (
    .a(al_ad19785e),
    .b(al_35a8bfef),
    .c(pause_source_addr[25]),
    .d(s_axi_wdata[25]),
    .e(al_868a1cad[25]),
    .o(al_238a702c[25]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_f9bda9db (
    .a(al_ad19785e),
    .b(al_35a8bfef),
    .c(pause_source_addr[26]),
    .d(s_axi_wdata[26]),
    .e(al_868a1cad[26]),
    .o(al_238a702c[26]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_db413542 (
    .a(al_ad19785e),
    .b(al_35a8bfef),
    .c(pause_source_addr[27]),
    .d(s_axi_wdata[27]),
    .e(al_868a1cad[27]),
    .o(al_238a702c[27]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_ada16de9 (
    .a(al_ad19785e),
    .b(al_35a8bfef),
    .c(pause_source_addr[28]),
    .d(s_axi_wdata[28]),
    .e(al_868a1cad[28]),
    .o(al_238a702c[28]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_3b39753 (
    .a(al_ad19785e),
    .b(al_35a8bfef),
    .c(pause_source_addr[29]),
    .d(s_axi_wdata[29]),
    .e(al_868a1cad[29]),
    .o(al_238a702c[29]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_6174330d (
    .a(al_ad19785e),
    .b(al_35a8bfef),
    .c(pause_source_addr[2]),
    .d(s_axi_wdata[2]),
    .e(al_868a1cad[2]),
    .o(al_238a702c[2]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*B*A)"),
    .INIT(32'h00000080))
    al_fa9a871c (
    .a(al_cf696ef0),
    .b(al_13660933[4]),
    .c(al_13660933[5]),
    .d(al_13660933[6]),
    .e(al_13660933[7]),
    .o(al_ad19785e));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_fcc6cbe (
    .a(al_ad19785e),
    .b(al_35a8bfef),
    .c(pause_source_addr[30]),
    .d(s_axi_wdata[30]),
    .e(al_868a1cad[30]),
    .o(al_238a702c[30]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_c370187d (
    .a(al_ad19785e),
    .b(al_35a8bfef),
    .c(pause_source_addr[31]),
    .d(s_axi_wdata[31]),
    .e(al_868a1cad[31]),
    .o(al_238a702c[31]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_982e9058 (
    .a(al_ad19785e),
    .b(al_35a8bfef),
    .c(pause_source_addr[3]),
    .d(s_axi_wdata[3]),
    .e(al_868a1cad[3]),
    .o(al_238a702c[3]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_cc5d6f6e (
    .a(al_ad19785e),
    .b(al_35a8bfef),
    .c(pause_source_addr[4]),
    .d(s_axi_wdata[4]),
    .e(al_868a1cad[4]),
    .o(al_238a702c[4]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_2c876d80 (
    .a(al_ad19785e),
    .b(al_35a8bfef),
    .c(pause_source_addr[5]),
    .d(s_axi_wdata[5]),
    .e(al_868a1cad[5]),
    .o(al_238a702c[5]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_aa233441 (
    .a(al_ad19785e),
    .b(al_35a8bfef),
    .c(pause_source_addr[6]),
    .d(s_axi_wdata[6]),
    .e(al_868a1cad[6]),
    .o(al_238a702c[6]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_7565903c (
    .a(al_ad19785e),
    .b(al_35a8bfef),
    .c(pause_source_addr[7]),
    .d(s_axi_wdata[7]),
    .e(al_868a1cad[7]),
    .o(al_238a702c[7]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_74783b59 (
    .a(al_ad19785e),
    .b(al_35a8bfef),
    .c(pause_source_addr[8]),
    .d(s_axi_wdata[8]),
    .e(al_868a1cad[8]),
    .o(al_238a702c[8]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_f7ab217b (
    .a(al_ad19785e),
    .b(al_35a8bfef),
    .c(pause_source_addr[9]),
    .d(s_axi_wdata[9]),
    .e(al_868a1cad[9]),
    .o(al_238a702c[9]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_4f3dd0b7 (
    .a(al_1c908f3d),
    .b(al_35a8bfef),
    .c(pause_source_addr[32]),
    .d(s_axi_wdata[0]),
    .e(al_cd0aa0ee[0]),
    .o(al_939ca227[0]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_c2eef666 (
    .a(al_1c908f3d),
    .b(al_35a8bfef),
    .c(pause_source_addr[42]),
    .d(s_axi_wdata[10]),
    .e(al_cd0aa0ee[10]),
    .o(al_939ca227[10]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_dd82c1c2 (
    .a(al_1c908f3d),
    .b(al_35a8bfef),
    .c(pause_source_addr[43]),
    .d(s_axi_wdata[11]),
    .e(al_cd0aa0ee[11]),
    .o(al_939ca227[11]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_40e3e1d8 (
    .a(al_1c908f3d),
    .b(al_35a8bfef),
    .c(pause_source_addr[44]),
    .d(s_axi_wdata[12]),
    .e(al_cd0aa0ee[12]),
    .o(al_939ca227[12]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_61efc3a (
    .a(al_1c908f3d),
    .b(al_35a8bfef),
    .c(pause_source_addr[45]),
    .d(s_axi_wdata[13]),
    .e(al_cd0aa0ee[13]),
    .o(al_939ca227[13]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_c00d79ec (
    .a(al_81344cef),
    .b(al_a0f12bef[0]),
    .o(al_35a8bfef));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*~C*~B*A)"),
    .INIT(32'h00000200))
    al_1d81858c (
    .a(al_cf696ef0),
    .b(al_13660933[4]),
    .c(al_13660933[5]),
    .d(al_13660933[6]),
    .e(al_13660933[7]),
    .o(al_1c908f3d));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_80ac601 (
    .a(al_1c908f3d),
    .b(al_35a8bfef),
    .c(pause_source_addr[46]),
    .d(s_axi_wdata[14]),
    .e(al_cd0aa0ee[14]),
    .o(al_939ca227[14]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_2548590 (
    .a(al_1c908f3d),
    .b(al_35a8bfef),
    .c(pause_source_addr[47]),
    .d(s_axi_wdata[15]),
    .e(al_cd0aa0ee[15]),
    .o(al_939ca227[15]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_8022701c (
    .a(al_1c908f3d),
    .b(al_35a8bfef),
    .c(pause_source_addr[33]),
    .d(s_axi_wdata[1]),
    .e(al_cd0aa0ee[1]),
    .o(al_939ca227[1]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_c2f29361 (
    .a(al_1c908f3d),
    .b(al_35a8bfef),
    .c(pause_source_addr[34]),
    .d(s_axi_wdata[2]),
    .e(al_cd0aa0ee[2]),
    .o(al_939ca227[2]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_f4cf8c4a (
    .a(al_1c908f3d),
    .b(al_35a8bfef),
    .c(pause_source_addr[35]),
    .d(s_axi_wdata[3]),
    .e(al_cd0aa0ee[3]),
    .o(al_939ca227[3]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_ec1f1435 (
    .a(al_1c908f3d),
    .b(al_35a8bfef),
    .c(pause_source_addr[36]),
    .d(s_axi_wdata[4]),
    .e(al_cd0aa0ee[4]),
    .o(al_939ca227[4]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_1094d0c0 (
    .a(al_1c908f3d),
    .b(al_35a8bfef),
    .c(pause_source_addr[37]),
    .d(s_axi_wdata[5]),
    .e(al_cd0aa0ee[5]),
    .o(al_939ca227[5]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_b7d677d2 (
    .a(al_1c908f3d),
    .b(al_35a8bfef),
    .c(pause_source_addr[38]),
    .d(s_axi_wdata[6]),
    .e(al_cd0aa0ee[6]),
    .o(al_939ca227[6]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_eed70f94 (
    .a(al_1c908f3d),
    .b(al_35a8bfef),
    .c(pause_source_addr[39]),
    .d(s_axi_wdata[7]),
    .e(al_cd0aa0ee[7]),
    .o(al_939ca227[7]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_88c24801 (
    .a(al_1c908f3d),
    .b(al_35a8bfef),
    .c(pause_source_addr[40]),
    .d(s_axi_wdata[8]),
    .e(al_cd0aa0ee[8]),
    .o(al_939ca227[8]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    al_1ace6dfd (
    .a(al_1c908f3d),
    .b(al_35a8bfef),
    .c(pause_source_addr[41]),
    .d(s_axi_wdata[9]),
    .e(al_cd0aa0ee[9]),
    .o(al_939ca227[9]));
  AL_MAP_LUT5 #(
    .EQN("(E*D*~C*~B*A)"),
    .INIT(32'h02000000))
    al_5f08a234 (
    .a(al_cf696ef0),
    .b(al_13660933[4]),
    .c(al_13660933[5]),
    .d(al_13660933[6]),
    .e(al_13660933[7]),
    .o(al_1ce50ae3));
  AL_MAP_LUT4 #(
    .EQN("((~D*C)*~(B)*~(A)+(~D*C)*B*~(A)+~((~D*C))*B*A+(~D*C)*B*A)"),
    .INIT(16'h88d8))
    al_5b9e417 (
    .a(al_dbd330f5),
    .b(s_axi_awaddr[0]),
    .c(al_13660933[0]),
    .d(s_axi_bvalid),
    .o(al_3833d624[0]));
  AL_MAP_LUT4 #(
    .EQN("((~D*C)*~(B)*~(A)+(~D*C)*B*~(A)+~((~D*C))*B*A+(~D*C)*B*A)"),
    .INIT(16'h88d8))
    al_7a9542a3 (
    .a(al_dbd330f5),
    .b(s_axi_awaddr[1]),
    .c(al_13660933[1]),
    .d(s_axi_bvalid),
    .o(al_3833d624[1]));
  AL_MAP_LUT4 #(
    .EQN("((~D*C)*~(B)*~(A)+(~D*C)*B*~(A)+~((~D*C))*B*A+(~D*C)*B*A)"),
    .INIT(16'h88d8))
    al_f8b8275 (
    .a(al_dbd330f5),
    .b(s_axi_awaddr[2]),
    .c(al_13660933[2]),
    .d(s_axi_bvalid),
    .o(al_3833d624[2]));
  AL_MAP_LUT4 #(
    .EQN("((~D*C)*~(B)*~(A)+(~D*C)*B*~(A)+~((~D*C))*B*A+(~D*C)*B*A)"),
    .INIT(16'h88d8))
    al_a9668d1b (
    .a(al_dbd330f5),
    .b(s_axi_awaddr[3]),
    .c(al_13660933[3]),
    .d(s_axi_bvalid),
    .o(al_3833d624[3]));
  AL_MAP_LUT4 #(
    .EQN("((~D*C)*~(B)*~(A)+(~D*C)*B*~(A)+~((~D*C))*B*A+(~D*C)*B*A)"),
    .INIT(16'h88d8))
    al_f0c236bd (
    .a(al_dbd330f5),
    .b(s_axi_awaddr[4]),
    .c(al_13660933[4]),
    .d(s_axi_bvalid),
    .o(al_3833d624[4]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_45f46f3c (
    .a(s_axi_awvalid),
    .b(s_axi_wvalid),
    .c(s_axi_wready),
    .o(al_dbd330f5));
  AL_MAP_LUT4 #(
    .EQN("((~D*C)*~(B)*~(A)+(~D*C)*B*~(A)+~((~D*C))*B*A+(~D*C)*B*A)"),
    .INIT(16'h88d8))
    al_36754613 (
    .a(al_dbd330f5),
    .b(s_axi_awaddr[5]),
    .c(al_13660933[5]),
    .d(s_axi_bvalid),
    .o(al_3833d624[5]));
  AL_MAP_LUT4 #(
    .EQN("((~D*C)*~(B)*~(A)+(~D*C)*B*~(A)+~((~D*C))*B*A+(~D*C)*B*A)"),
    .INIT(16'h88d8))
    al_d95ab129 (
    .a(al_dbd330f5),
    .b(s_axi_awaddr[6]),
    .c(al_13660933[6]),
    .d(s_axi_bvalid),
    .o(al_3833d624[6]));
  AL_MAP_LUT4 #(
    .EQN("((~D*C)*~(B)*~(A)+(~D*C)*B*~(A)+~((~D*C))*B*A+(~D*C)*B*A)"),
    .INIT(16'h88d8))
    al_16e13987 (
    .a(al_dbd330f5),
    .b(s_axi_awaddr[7]),
    .c(al_13660933[7]),
    .d(s_axi_bvalid),
    .o(al_3833d624[7]));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*B*~(C)*~(D)*~((F*~E))+~(A)*B*C*~(D)*~((F*~E))+~(A)*~(B)*~(C)*D*~((F*~E))+A*~(B)*~(C)*D*~((F*~E))+~(A)*B*~(C)*D*~((F*~E))+A*B*~(C)*D*~((F*~E))+A*~(B)*~(C)*~(D)*(F*~E)+~(A)*B*~(C)*~(D)*(F*~E)+A*B*~(C)*~(D)*(F*~E)+A*~(B)*C*~(D)*(F*~E)+~(A)*B*C*~(D)*(F*~E)+A*B*C*~(D)*(F*~E)+~(A)*~(B)*~(C)*D*(F*~E)+A*~(B)*~(C)*D*(F*~E)+~(A)*B*~(C)*D*(F*~E)+A*B*~(C)*D*(F*~E)+A*~(B)*C*D*(F*~E)+A*B*C*D*(F*~E))"),
    .INIT(64'h0f44afee0f440f44))
    al_458b0ece (
    .a(al_5d31465b),
    .b(al_5df5c44f),
    .c(s_axi_bready),
    .d(s_axi_bvalid),
    .e(al_2b48f483),
    .f(al_841146bf),
    .o(al_bf676c3e));
  AL_MAP_LUT4 #(
    .EQN("((~D*C)*~(B)*~(A)+(~D*C)*B*~(A)+~((~D*C))*B*A+(~D*C)*B*A)"),
    .INIT(16'h88d8))
    al_94ead4d1 (
    .a(al_a584e1fd),
    .b(s_axi_araddr[0]),
    .c(al_82716c38[0]),
    .d(s_axi_rvalid),
    .o(al_7b2ceef0[0]));
  AL_MAP_LUT4 #(
    .EQN("((~D*C)*~(B)*~(A)+(~D*C)*B*~(A)+~((~D*C))*B*A+(~D*C)*B*A)"),
    .INIT(16'h88d8))
    al_ee60e615 (
    .a(al_a584e1fd),
    .b(s_axi_araddr[1]),
    .c(al_82716c38[1]),
    .d(s_axi_rvalid),
    .o(al_7b2ceef0[1]));
  AL_MAP_LUT4 #(
    .EQN("((~D*C)*~(B)*~(A)+(~D*C)*B*~(A)+~((~D*C))*B*A+(~D*C)*B*A)"),
    .INIT(16'h88d8))
    al_c496b1da (
    .a(al_a584e1fd),
    .b(s_axi_araddr[2]),
    .c(al_82716c38[2]),
    .d(s_axi_rvalid),
    .o(al_7b2ceef0[2]));
  AL_MAP_LUT4 #(
    .EQN("((~D*C)*~(B)*~(A)+(~D*C)*B*~(A)+~((~D*C))*B*A+(~D*C)*B*A)"),
    .INIT(16'h88d8))
    al_d3311b4e (
    .a(al_a584e1fd),
    .b(s_axi_araddr[3]),
    .c(al_82716c38[3]),
    .d(s_axi_rvalid),
    .o(al_7b2ceef0[3]));
  AL_MAP_LUT4 #(
    .EQN("((~D*C)*~(B)*~(A)+(~D*C)*B*~(A)+~((~D*C))*B*A+(~D*C)*B*A)"),
    .INIT(16'h88d8))
    al_6ea7427d (
    .a(al_a584e1fd),
    .b(s_axi_araddr[4]),
    .c(al_82716c38[4]),
    .d(s_axi_rvalid),
    .o(al_7b2ceef0[4]));
  AL_MAP_LUT4 #(
    .EQN("((~D*C)*~(B)*~(A)+(~D*C)*B*~(A)+~((~D*C))*B*A+(~D*C)*B*A)"),
    .INIT(16'h88d8))
    al_5756b039 (
    .a(al_a584e1fd),
    .b(s_axi_araddr[5]),
    .c(al_82716c38[5]),
    .d(s_axi_rvalid),
    .o(al_7b2ceef0[5]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_53eabc02 (
    .a(s_axi_arvalid),
    .b(s_axi_arready),
    .o(al_a584e1fd));
  AL_MAP_LUT4 #(
    .EQN("((~D*C)*~(B)*~(A)+(~D*C)*B*~(A)+~((~D*C))*B*A+(~D*C)*B*A)"),
    .INIT(16'h88d8))
    al_8e517a73 (
    .a(al_a584e1fd),
    .b(s_axi_araddr[6]),
    .c(al_82716c38[6]),
    .d(s_axi_rvalid),
    .o(al_7b2ceef0[6]));
  AL_MAP_LUT4 #(
    .EQN("((~D*C)*~(B)*~(A)+(~D*C)*B*~(A)+~((~D*C))*B*A+(~D*C)*B*A)"),
    .INIT(16'h88d8))
    al_9ac71553 (
    .a(al_a584e1fd),
    .b(s_axi_araddr[7]),
    .c(al_82716c38[7]),
    .d(s_axi_rvalid),
    .o(al_7b2ceef0[7]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_e2c8c09c (
    .a(s_axi_arvalid),
    .b(s_axi_arready),
    .c(s_axi_rvalid),
    .o(al_e8564782));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*C*~B*A)"),
    .INIT(32'h00200000))
    al_879ec194 (
    .a(al_711bc49b),
    .b(al_82716c38[4]),
    .c(al_82716c38[5]),
    .d(al_82716c38[6]),
    .e(al_82716c38[7]),
    .o(al_2086b792));
  AL_MAP_LUT6 #(
    .EQN("~(~(D*~C)*~(B*~((F*~E))*~(A)+B*(F*~E)*~(A)+~(B)*(F*~E)*A+B*(F*~E)*A))"),
    .INIT(64'h4f44efee4f444f44))
    al_4490efaf (
    .a(al_2086b792),
    .b(al_e8564782),
    .c(s_axi_rready),
    .d(s_axi_rvalid),
    .e(al_2b48f483),
    .f(al_841146bf),
    .o(al_1d703c48));
  AL_DFF_X al_a209e4a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_82626899),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a9406400));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*C*B*A)"),
    .INIT(32'h00008000))
    al_15f26e6d (
    .a(al_cf696ef0),
    .b(al_13660933[4]),
    .c(al_13660933[5]),
    .d(al_13660933[6]),
    .e(al_13660933[7]),
    .o(al_57e16e6f));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'hfdf8))
    al_30685efe (
    .a(al_57e16e6f),
    .b(s_axi_wdata[0]),
    .c(al_81344cef),
    .d(al_a9406400),
    .o(al_82626899));
  AL_DFF_X al_dacd13c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_3833d624[0]),
    .en(1'b1),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_13660933[0]));
  AL_DFF_X al_46a68ad8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_3833d624[1]),
    .en(1'b1),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_13660933[1]));
  AL_DFF_X al_63682572 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_3833d624[2]),
    .en(1'b1),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_13660933[2]));
  AL_DFF_X al_1d022814 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_3833d624[3]),
    .en(1'b1),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_13660933[3]));
  AL_DFF_X al_bee0e0d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_3833d624[4]),
    .en(1'b1),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_13660933[4]));
  AL_DFF_X al_b2f0bc26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_3833d624[5]),
    .en(1'b1),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_13660933[5]));
  AL_DFF_X al_866dd369 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_3833d624[6]),
    .en(1'b1),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_13660933[6]));
  AL_DFF_X al_5d44bc9c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_3833d624[7]),
    .en(1'b1),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_13660933[7]));
  AL_DFF_X al_554b625 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_7b2ceef0[0]),
    .en(1'b1),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_82716c38[0]));
  AL_DFF_X al_358b1dce (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_7b2ceef0[1]),
    .en(1'b1),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_82716c38[1]));
  AL_DFF_X al_d7cebac8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_7b2ceef0[2]),
    .en(1'b1),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_82716c38[2]));
  AL_DFF_X al_d2ce4dcf (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_7b2ceef0[3]),
    .en(1'b1),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_82716c38[3]));
  AL_DFF_X al_32b6d60b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_7b2ceef0[4]),
    .en(1'b1),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_82716c38[4]));
  AL_DFF_X al_ba6b982f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_7b2ceef0[5]),
    .en(1'b1),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_82716c38[5]));
  AL_DFF_X al_e91bead3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_7b2ceef0[6]),
    .en(1'b1),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_82716c38[6]));
  AL_DFF_X al_48b59abf (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_7b2ceef0[7]),
    .en(1'b1),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_82716c38[7]));
  AL_DFF_X al_a3c3c524 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_492d1bb8[0]),
    .en(al_e8564782),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_88fb5330[0]));
  AL_DFF_X al_99c65a0e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_492d1bb8[9]),
    .en(al_e8564782),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_88fb5330[9]));
  AL_DFF_X al_d165124d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_492d1bb8[10]),
    .en(al_e8564782),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_88fb5330[10]));
  AL_DFF_X al_287a92ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_492d1bb8[11]),
    .en(al_e8564782),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_88fb5330[11]));
  AL_DFF_X al_a76d0050 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_492d1bb8[12]),
    .en(al_e8564782),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_88fb5330[12]));
  AL_DFF_X al_db2f7aab (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_492d1bb8[13]),
    .en(al_e8564782),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_88fb5330[13]));
  AL_DFF_X al_45f13ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_492d1bb8[14]),
    .en(al_e8564782),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_88fb5330[14]));
  AL_DFF_X al_b1228db6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_492d1bb8[15]),
    .en(al_e8564782),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_88fb5330[15]));
  AL_DFF_X al_83dba831 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_492d1bb8[16]),
    .en(al_e8564782),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_88fb5330[16]));
  AL_DFF_X al_40a38860 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_492d1bb8[17]),
    .en(al_e8564782),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_88fb5330[17]));
  AL_DFF_X al_a1d35d32 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_492d1bb8[18]),
    .en(al_e8564782),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_88fb5330[18]));
  AL_DFF_X al_b7e4b655 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_492d1bb8[1]),
    .en(al_e8564782),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_88fb5330[1]));
  AL_DFF_X al_1d12639a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_492d1bb8[19]),
    .en(al_e8564782),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_88fb5330[19]));
  AL_DFF_X al_32d7a679 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_492d1bb8[20]),
    .en(al_e8564782),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_88fb5330[20]));
  AL_DFF_X al_8ac1f791 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_492d1bb8[21]),
    .en(al_e8564782),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_88fb5330[21]));
  AL_DFF_X al_27ab96d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_492d1bb8[22]),
    .en(al_e8564782),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_88fb5330[22]));
  AL_DFF_X al_fa81d69 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_492d1bb8[23]),
    .en(al_e8564782),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_88fb5330[23]));
  AL_DFF_X al_3c4ef7ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_492d1bb8[24]),
    .en(al_e8564782),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_88fb5330[24]));
  AL_DFF_X al_f3ed6b2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_492d1bb8[25]),
    .en(al_e8564782),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_88fb5330[25]));
  AL_DFF_X al_7ecd582c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_492d1bb8[26]),
    .en(al_e8564782),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_88fb5330[26]));
  AL_DFF_X al_65ca0477 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_492d1bb8[27]),
    .en(al_e8564782),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_88fb5330[27]));
  AL_DFF_X al_89d557a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_492d1bb8[28]),
    .en(al_e8564782),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_88fb5330[28]));
  AL_DFF_X al_2c4c4eeb (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_492d1bb8[2]),
    .en(al_e8564782),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_88fb5330[2]));
  AL_DFF_X al_2bb485ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_492d1bb8[29]),
    .en(al_e8564782),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_88fb5330[29]));
  AL_DFF_X al_157363e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_492d1bb8[30]),
    .en(al_e8564782),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_88fb5330[30]));
  AL_DFF_X al_ca0b60d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_492d1bb8[31]),
    .en(al_e8564782),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_88fb5330[31]));
  AL_DFF_X al_8f85979d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_492d1bb8[3]),
    .en(al_e8564782),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_88fb5330[3]));
  AL_DFF_X al_95f7d71e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_492d1bb8[4]),
    .en(al_e8564782),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_88fb5330[4]));
  AL_DFF_X al_8f4456c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_492d1bb8[5]),
    .en(al_e8564782),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_88fb5330[5]));
  AL_DFF_X al_ee3f784f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_492d1bb8[6]),
    .en(al_e8564782),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_88fb5330[6]));
  AL_DFF_X al_86681e08 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_492d1bb8[7]),
    .en(al_e8564782),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_88fb5330[7]));
  AL_DFF_X al_4be618f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_492d1bb8[8]),
    .en(al_e8564782),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_88fb5330[8]));
  AL_DFF_X al_9511645c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_e7647890),
    .en(1'b1),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_9b4eaefc[0]));
  AL_DFF_X al_5de664dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[9]),
    .en(al_c3d9ce92),
    .sr(al_1b655917),
    .ss(1'b0),
    .q(al_9b4eaefc[9]));
  AL_DFF_X al_3145d5b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[10]),
    .en(al_c3d9ce92),
    .sr(al_1b655917),
    .ss(1'b0),
    .q(al_9b4eaefc[10]));
  AL_DFF_X al_dd8d06f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[11]),
    .en(al_c3d9ce92),
    .sr(al_1b655917),
    .ss(1'b0),
    .q(al_9b4eaefc[11]));
  AL_DFF_X al_769e813c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[12]),
    .en(al_c3d9ce92),
    .sr(al_1b655917),
    .ss(1'b0),
    .q(al_9b4eaefc[12]));
  AL_DFF_X al_d4de155a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[13]),
    .en(al_c3d9ce92),
    .sr(al_1b655917),
    .ss(1'b0),
    .q(al_9b4eaefc[13]));
  AL_DFF_X al_c1f42121 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[14]),
    .en(al_c3d9ce92),
    .sr(al_1b655917),
    .ss(1'b0),
    .q(al_9b4eaefc[14]));
  AL_DFF_X al_cb24c1b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[15]),
    .en(al_c3d9ce92),
    .sr(al_1b655917),
    .ss(1'b0),
    .q(al_9b4eaefc[15]));
  AL_DFF_X al_990fc3de (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[16]),
    .en(al_c3d9ce92),
    .sr(al_1b655917),
    .ss(1'b0),
    .q(al_9b4eaefc[16]));
  AL_DFF_X al_82de513 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[17]),
    .en(al_c3d9ce92),
    .sr(al_1b655917),
    .ss(1'b0),
    .q(al_9b4eaefc[17]));
  AL_DFF_X al_3825819c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[18]),
    .en(al_c3d9ce92),
    .sr(al_1b655917),
    .ss(1'b0),
    .q(al_9b4eaefc[18]));
  AL_DFF_X al_b0c360af (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[1]),
    .en(al_c3d9ce92),
    .sr(1'b0),
    .ss(al_1b655917),
    .q(al_9b4eaefc[1]));
  AL_DFF_X al_ea24b8ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[19]),
    .en(al_c3d9ce92),
    .sr(al_1b655917),
    .ss(1'b0),
    .q(al_9b4eaefc[19]));
  AL_DFF_X al_81d929ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[20]),
    .en(al_c3d9ce92),
    .sr(al_1b655917),
    .ss(1'b0),
    .q(al_9b4eaefc[20]));
  AL_DFF_X al_9556d7db (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[21]),
    .en(al_c3d9ce92),
    .sr(al_1b655917),
    .ss(1'b0),
    .q(al_9b4eaefc[21]));
  AL_DFF_X al_cc2a365f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[22]),
    .en(al_c3d9ce92),
    .sr(al_1b655917),
    .ss(1'b0),
    .q(al_9b4eaefc[22]));
  AL_DFF_X al_4a79c48b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[23]),
    .en(al_c3d9ce92),
    .sr(al_1b655917),
    .ss(1'b0),
    .q(al_9b4eaefc[23]));
  AL_DFF_X al_e1b20d2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[24]),
    .en(al_c3d9ce92),
    .sr(al_1b655917),
    .ss(1'b0),
    .q(al_9b4eaefc[24]));
  AL_DFF_X al_cf28748d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[25]),
    .en(al_c3d9ce92),
    .sr(al_1b655917),
    .ss(1'b0),
    .q(al_9b4eaefc[25]));
  AL_DFF_X al_69db6114 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[26]),
    .en(al_c3d9ce92),
    .sr(al_1b655917),
    .ss(1'b0),
    .q(al_9b4eaefc[26]));
  AL_DFF_X al_ea79fbe0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[27]),
    .en(al_c3d9ce92),
    .sr(al_1b655917),
    .ss(1'b0),
    .q(al_9b4eaefc[27]));
  AL_DFF_X al_2eaadbe6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[28]),
    .en(al_c3d9ce92),
    .sr(al_1b655917),
    .ss(1'b0),
    .q(al_9b4eaefc[28]));
  AL_DFF_X al_b884dfe7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[2]),
    .en(al_c3d9ce92),
    .sr(al_1b655917),
    .ss(1'b0),
    .q(al_9b4eaefc[2]));
  AL_DFF_X al_f1629e2c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[29]),
    .en(al_c3d9ce92),
    .sr(al_1b655917),
    .ss(1'b0),
    .q(al_9b4eaefc[29]));
  AL_DFF_X al_e5397a0c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[30]),
    .en(al_c3d9ce92),
    .sr(al_1b655917),
    .ss(1'b0),
    .q(al_9b4eaefc[30]));
  AL_DFF_X al_1ea68e95 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[31]),
    .en(al_c3d9ce92),
    .sr(al_1b655917),
    .ss(1'b0),
    .q(al_9b4eaefc[31]));
  AL_DFF_X al_18e0716d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[3]),
    .en(al_c3d9ce92),
    .sr(al_1b655917),
    .ss(1'b0),
    .q(al_9b4eaefc[3]));
  AL_DFF_X al_3ead7d8a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[4]),
    .en(al_c3d9ce92),
    .sr(al_1b655917),
    .ss(1'b0),
    .q(al_9b4eaefc[4]));
  AL_DFF_X al_43088097 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[5]),
    .en(al_c3d9ce92),
    .sr(al_1b655917),
    .ss(1'b0),
    .q(al_9b4eaefc[5]));
  AL_DFF_X al_5172ac84 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[6]),
    .en(al_c3d9ce92),
    .sr(al_1b655917),
    .ss(1'b0),
    .q(al_9b4eaefc[6]));
  AL_DFF_X al_965c0b5d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[7]),
    .en(al_c3d9ce92),
    .sr(al_1b655917),
    .ss(1'b0),
    .q(al_9b4eaefc[7]));
  AL_DFF_X al_ad73dfca (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[8]),
    .en(al_c3d9ce92),
    .sr(al_1b655917),
    .ss(1'b0),
    .q(al_9b4eaefc[8]));
  AL_DFF_X al_79656483 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_624c8b6f),
    .en(1'b1),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_a0f12bef[0]));
  AL_DFF_X al_b5ddf65f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[9]),
    .en(al_291f5813),
    .sr(al_35a8bfef),
    .ss(1'b0),
    .q(al_a0f12bef[9]));
  AL_DFF_X al_daf0bc3f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[10]),
    .en(al_291f5813),
    .sr(al_35a8bfef),
    .ss(1'b0),
    .q(al_a0f12bef[10]));
  AL_DFF_X al_ce546bd3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[11]),
    .en(al_291f5813),
    .sr(al_35a8bfef),
    .ss(1'b0),
    .q(al_a0f12bef[11]));
  AL_DFF_X al_5f4bb1fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[12]),
    .en(al_291f5813),
    .sr(al_35a8bfef),
    .ss(1'b0),
    .q(al_a0f12bef[12]));
  AL_DFF_X al_f69fa14d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[13]),
    .en(al_291f5813),
    .sr(al_35a8bfef),
    .ss(1'b0),
    .q(al_a0f12bef[13]));
  AL_DFF_X al_cf45c72e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[14]),
    .en(al_291f5813),
    .sr(al_35a8bfef),
    .ss(1'b0),
    .q(al_a0f12bef[14]));
  AL_DFF_X al_a631d4fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[15]),
    .en(al_291f5813),
    .sr(al_35a8bfef),
    .ss(1'b0),
    .q(al_a0f12bef[15]));
  AL_DFF_X al_560b110c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[16]),
    .en(al_291f5813),
    .sr(al_35a8bfef),
    .ss(1'b0),
    .q(al_a0f12bef[16]));
  AL_DFF_X al_92415293 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[17]),
    .en(al_291f5813),
    .sr(al_35a8bfef),
    .ss(1'b0),
    .q(al_a0f12bef[17]));
  AL_DFF_X al_6cce0f4a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[18]),
    .en(al_291f5813),
    .sr(al_35a8bfef),
    .ss(1'b0),
    .q(al_a0f12bef[18]));
  AL_DFF_X al_ee82d183 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[1]),
    .en(al_291f5813),
    .sr(1'b0),
    .ss(al_35a8bfef),
    .q(al_a0f12bef[1]));
  AL_DFF_X al_2caa66e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[19]),
    .en(al_291f5813),
    .sr(al_35a8bfef),
    .ss(1'b0),
    .q(al_a0f12bef[19]));
  AL_DFF_X al_73594816 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[20]),
    .en(al_291f5813),
    .sr(al_35a8bfef),
    .ss(1'b0),
    .q(al_a0f12bef[20]));
  AL_DFF_X al_bf5bcb1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[21]),
    .en(al_291f5813),
    .sr(al_35a8bfef),
    .ss(1'b0),
    .q(al_a0f12bef[21]));
  AL_DFF_X al_cb6594aa (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[22]),
    .en(al_291f5813),
    .sr(al_35a8bfef),
    .ss(1'b0),
    .q(al_a0f12bef[22]));
  AL_DFF_X al_9d074962 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[23]),
    .en(al_291f5813),
    .sr(al_35a8bfef),
    .ss(1'b0),
    .q(al_a0f12bef[23]));
  AL_DFF_X al_12998340 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[24]),
    .en(al_291f5813),
    .sr(al_35a8bfef),
    .ss(1'b0),
    .q(al_a0f12bef[24]));
  AL_DFF_X al_8de1afac (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[25]),
    .en(al_291f5813),
    .sr(al_35a8bfef),
    .ss(1'b0),
    .q(al_a0f12bef[25]));
  AL_DFF_X al_6b9c6db2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[26]),
    .en(al_291f5813),
    .sr(al_35a8bfef),
    .ss(1'b0),
    .q(al_a0f12bef[26]));
  AL_DFF_X al_9d039895 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[27]),
    .en(al_291f5813),
    .sr(al_35a8bfef),
    .ss(1'b0),
    .q(al_a0f12bef[27]));
  AL_DFF_X al_24e92dce (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[28]),
    .en(al_291f5813),
    .sr(al_35a8bfef),
    .ss(1'b0),
    .q(al_a0f12bef[28]));
  AL_DFF_X al_a08dab40 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[2]),
    .en(al_291f5813),
    .sr(al_35a8bfef),
    .ss(1'b0),
    .q(al_a0f12bef[2]));
  AL_DFF_X al_6ed3b5a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[29]),
    .en(al_291f5813),
    .sr(al_35a8bfef),
    .ss(1'b0),
    .q(al_a0f12bef[29]));
  AL_DFF_X al_5a4c4ebc (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[30]),
    .en(al_291f5813),
    .sr(al_35a8bfef),
    .ss(1'b0),
    .q(al_a0f12bef[30]));
  AL_DFF_X al_b1faf88 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[31]),
    .en(al_291f5813),
    .sr(al_35a8bfef),
    .ss(1'b0),
    .q(al_a0f12bef[31]));
  AL_DFF_X al_a066e66 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[3]),
    .en(al_291f5813),
    .sr(al_35a8bfef),
    .ss(1'b0),
    .q(al_a0f12bef[3]));
  AL_DFF_X al_ba794bb7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[4]),
    .en(al_291f5813),
    .sr(al_35a8bfef),
    .ss(1'b0),
    .q(al_a0f12bef[4]));
  AL_DFF_X al_d5d921c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[5]),
    .en(al_291f5813),
    .sr(al_35a8bfef),
    .ss(1'b0),
    .q(al_a0f12bef[5]));
  AL_DFF_X al_6eec50c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[6]),
    .en(al_291f5813),
    .sr(al_35a8bfef),
    .ss(1'b0),
    .q(al_a0f12bef[6]));
  AL_DFF_X al_ffe975a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[7]),
    .en(al_291f5813),
    .sr(al_35a8bfef),
    .ss(1'b0),
    .q(al_a0f12bef[7]));
  AL_DFF_X al_ebb40327 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[8]),
    .en(al_291f5813),
    .sr(al_35a8bfef),
    .ss(1'b0),
    .q(al_a0f12bef[8]));
  AL_DFF_X al_9972f7c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_238a702c[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_868a1cad[0]));
  AL_DFF_X al_528be1ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_238a702c[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_868a1cad[9]));
  AL_DFF_X al_33839558 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_238a702c[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_868a1cad[10]));
  AL_DFF_X al_35f62c44 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_238a702c[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_868a1cad[11]));
  AL_DFF_X al_34887c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_238a702c[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_868a1cad[12]));
  AL_DFF_X al_5100591c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_238a702c[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_868a1cad[13]));
  AL_DFF_X al_c54785f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_238a702c[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_868a1cad[14]));
  AL_DFF_X al_b2bf06c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_238a702c[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_868a1cad[15]));
  AL_DFF_X al_1a448de4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_238a702c[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_868a1cad[16]));
  AL_DFF_X al_3f671b60 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_238a702c[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_868a1cad[17]));
  AL_DFF_X al_db52d76d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_238a702c[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_868a1cad[18]));
  AL_DFF_X al_977fbc85 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_238a702c[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_868a1cad[1]));
  AL_DFF_X al_69f09ee0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_238a702c[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_868a1cad[19]));
  AL_DFF_X al_517921f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_238a702c[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_868a1cad[20]));
  AL_DFF_X al_d0aeeec0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_238a702c[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_868a1cad[21]));
  AL_DFF_X al_4479a350 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_238a702c[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_868a1cad[22]));
  AL_DFF_X al_f91d6ec6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_238a702c[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_868a1cad[23]));
  AL_DFF_X al_ad04bbe0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_238a702c[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_868a1cad[24]));
  AL_DFF_X al_1f7e4d44 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_238a702c[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_868a1cad[25]));
  AL_DFF_X al_f021522b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_238a702c[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_868a1cad[26]));
  AL_DFF_X al_c8cda48 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_238a702c[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_868a1cad[27]));
  AL_DFF_X al_3c4ff597 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_238a702c[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_868a1cad[28]));
  AL_DFF_X al_f71dbb93 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_238a702c[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_868a1cad[2]));
  AL_DFF_X al_841ebb0f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_238a702c[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_868a1cad[29]));
  AL_DFF_X al_7989aef4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_238a702c[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_868a1cad[30]));
  AL_DFF_X al_d091317d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_238a702c[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_868a1cad[31]));
  AL_DFF_X al_b9096d88 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_238a702c[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_868a1cad[3]));
  AL_DFF_X al_adffd074 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_238a702c[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_868a1cad[4]));
  AL_DFF_X al_9a1c2c9f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_238a702c[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_868a1cad[5]));
  AL_DFF_X al_2d71d89b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_238a702c[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_868a1cad[6]));
  AL_DFF_X al_744a0366 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_238a702c[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_868a1cad[7]));
  AL_DFF_X al_49cd3853 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_238a702c[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_868a1cad[8]));
  AL_DFF_X al_79a7d9bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_939ca227[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd0aa0ee[0]));
  AL_DFF_X al_26f57eec (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_939ca227[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd0aa0ee[9]));
  AL_DFF_X al_9f92ae4a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_939ca227[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd0aa0ee[10]));
  AL_DFF_X al_79effd38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_939ca227[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd0aa0ee[11]));
  AL_DFF_X al_53765b68 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_939ca227[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd0aa0ee[12]));
  AL_DFF_X al_216eb0c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_939ca227[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd0aa0ee[13]));
  AL_DFF_X al_a9b2139f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_939ca227[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd0aa0ee[14]));
  AL_DFF_X al_4eb4270a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_939ca227[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd0aa0ee[15]));
  AL_DFF_X al_c4d3b150 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_939ca227[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd0aa0ee[1]));
  AL_DFF_X al_8f568dea (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_939ca227[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd0aa0ee[2]));
  AL_DFF_X al_2da28edf (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_939ca227[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd0aa0ee[3]));
  AL_DFF_X al_7e50db2e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_939ca227[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd0aa0ee[4]));
  AL_DFF_X al_88479f6b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_939ca227[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd0aa0ee[5]));
  AL_DFF_X al_7a035f91 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_939ca227[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd0aa0ee[6]));
  AL_DFF_X al_d8deb4ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_939ca227[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd0aa0ee[7]));
  AL_DFF_X al_83e0a1e1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_939ca227[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cd0aa0ee[8]));
  AL_DFF_X al_4adb3463 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_43c0413c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25215c55[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_157b3e19 (
    .a(al_fc6dfd0c),
    .b(s_axi_wdata[1]),
    .c(al_25215c55[1]),
    .o(al_d94de5f0));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_f82f91 (
    .a(al_fc6dfd0c),
    .b(s_axi_wdata[0]),
    .c(al_25215c55[0]),
    .o(al_43c0413c));
  AL_DFF_X al_4a5ad6fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_d94de5f0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_25215c55[1]));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*~C*B*A)"),
    .INIT(32'h00000800))
    al_c074d5a4 (
    .a(al_cf696ef0),
    .b(al_13660933[4]),
    .c(al_13660933[5]),
    .d(al_13660933[6]),
    .e(al_13660933[7]),
    .o(al_fc6dfd0c));
  AL_DFF_X al_485a0b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_8f504dd9),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7808e039[0]));
  AL_DFF_X al_5aa06b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_7bf90fef),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7808e039[1]));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*C*~B*A)"),
    .INIT(32'h00002000))
    al_52107b89 (
    .a(al_cf696ef0),
    .b(al_13660933[4]),
    .c(al_13660933[5]),
    .d(al_13660933[6]),
    .e(al_13660933[7]),
    .o(al_2e19f5ba));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'hfdf8))
    al_59ffda02 (
    .a(al_2e19f5ba),
    .b(s_axi_wdata[0]),
    .c(al_81344cef),
    .d(al_7808e039[0]),
    .o(al_8f504dd9));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'hfdf8))
    al_4ffaadf1 (
    .a(al_2e19f5ba),
    .b(s_axi_wdata[1]),
    .c(al_81344cef),
    .d(al_7808e039[1]),
    .o(al_7bf90fef));
  AL_DFF_X al_5ee9dd42 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ec8f4956),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4096d0c7[0]));
  AL_DFF_X al_ee33bb06 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_d7d4dbcb),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4096d0c7[1]));
  AL_DFF_X al_e459b75c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_a97b8529),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4096d0c7[2]));
  AL_DFF_X al_b55ecd13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_dc2d168e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4096d0c7[3]));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    al_80ab4b9f (
    .a(al_cf696ef0),
    .b(al_41ffdcd4),
    .c(al_13660933[4]),
    .d(al_13660933[5]),
    .o(al_d5f82e51));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'h0d08))
    al_f1771e9c (
    .a(al_d5f82e51),
    .b(s_axi_wdata[0]),
    .c(al_81344cef),
    .d(al_4096d0c7[0]),
    .o(al_ec8f4956));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'hfdf8))
    al_fa2b99c7 (
    .a(al_d5f82e51),
    .b(s_axi_wdata[6]),
    .c(al_81344cef),
    .d(al_4096d0c7[6]),
    .o(al_495ff86c));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'h0d08))
    al_8a05bdef (
    .a(al_d5f82e51),
    .b(s_axi_wdata[5]),
    .c(al_81344cef),
    .d(al_4096d0c7[5]),
    .o(al_6dcc3ceb));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'h0d08))
    al_de6f0997 (
    .a(al_d5f82e51),
    .b(s_axi_wdata[4]),
    .c(al_81344cef),
    .d(al_4096d0c7[4]),
    .o(al_8127333f));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'h0d08))
    al_43e83449 (
    .a(al_d5f82e51),
    .b(s_axi_wdata[3]),
    .c(al_81344cef),
    .d(al_4096d0c7[3]),
    .o(al_dc2d168e));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'h0d08))
    al_c8113230 (
    .a(al_d5f82e51),
    .b(s_axi_wdata[2]),
    .c(al_81344cef),
    .d(al_4096d0c7[2]),
    .o(al_a97b8529));
  AL_DFF_X al_7f36a001 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_8127333f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4096d0c7[4]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'h0d08))
    al_29134af0 (
    .a(al_d5f82e51),
    .b(s_axi_wdata[1]),
    .c(al_81344cef),
    .d(al_4096d0c7[1]),
    .o(al_d7d4dbcb));
  AL_DFF_X al_6d437ae2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_6dcc3ceb),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4096d0c7[5]));
  AL_DFF_X al_976f0705 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_495ff86c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4096d0c7[6]));
  AL_DFF_X al_d76513f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_7a7f52dd),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_523025ae[0]));
  AL_DFF_X al_e8b9f205 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[9]),
    .en(al_3fec348f),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_523025ae[9]));
  AL_DFF_X al_ae303b67 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[10]),
    .en(al_3fec348f),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_523025ae[10]));
  AL_DFF_X al_3fd6996 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[11]),
    .en(al_3fec348f),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_523025ae[11]));
  AL_DFF_X al_7bf3518a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[12]),
    .en(al_3fec348f),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_523025ae[12]));
  AL_DFF_X al_c4188c82 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[1]),
    .en(al_3fec348f),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_523025ae[1]));
  AL_DFF_X al_806a6559 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[2]),
    .en(al_3fec348f),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_523025ae[2]));
  AL_DFF_X al_88c572fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[3]),
    .en(al_3fec348f),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_523025ae[3]));
  AL_DFF_X al_59875e34 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[4]),
    .en(al_3fec348f),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_523025ae[4]));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    al_147dcbbd (
    .a(al_13660933[2]),
    .b(al_13660933[3]),
    .c(al_13660933[4]),
    .d(al_13660933[5]),
    .o(al_a29e073));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_832639e6 (
    .a(al_a29e073),
    .b(al_41ffdcd4),
    .c(al_13660933[0]),
    .d(al_13660933[1]),
    .o(al_5d31465b));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_979c99bf (
    .a(al_5d31465b),
    .b(al_5df5c44f),
    .o(al_3fec348f));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_6dc17ca9 (
    .a(al_3fec348f),
    .b(s_axi_wdata[0]),
    .c(al_81344cef),
    .d(al_523025ae[0]),
    .o(al_7a7f52dd));
  AL_DFF_X al_c8a885f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[5]),
    .en(al_3fec348f),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_523025ae[5]));
  AL_DFF_X al_4dddfffa (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[6]),
    .en(al_3fec348f),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_523025ae[6]));
  AL_DFF_X al_cbdea2a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[7]),
    .en(al_3fec348f),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_523025ae[7]));
  AL_DFF_X al_a2cc2e1c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[8]),
    .en(al_3fec348f),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_523025ae[8]));
  AL_DFF_X al_7ab54f34 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[0]),
    .en(al_1ce50ae3),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_ab2a7f1[0]));
  AL_DFF_X al_d780dcf9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[9]),
    .en(al_1ce50ae3),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_ab2a7f1[9]));
  AL_DFF_X al_8317fddd (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[10]),
    .en(al_1ce50ae3),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_ab2a7f1[10]));
  AL_DFF_X al_88abef1a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[11]),
    .en(al_1ce50ae3),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_ab2a7f1[11]));
  AL_DFF_X al_f9d65d2f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[12]),
    .en(al_1ce50ae3),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_ab2a7f1[12]));
  AL_DFF_X al_e0310e1c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[13]),
    .en(al_1ce50ae3),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_ab2a7f1[13]));
  AL_DFF_X al_ddaff75b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[14]),
    .en(al_1ce50ae3),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_ab2a7f1[14]));
  AL_DFF_X al_a11d4d3b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[15]),
    .en(al_1ce50ae3),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_ab2a7f1[15]));
  AL_DFF_X al_15d17fb9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[1]),
    .en(al_1ce50ae3),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_ab2a7f1[1]));
  AL_DFF_X al_46fbf6c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[2]),
    .en(al_1ce50ae3),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_ab2a7f1[2]));
  AL_DFF_X al_1bc98316 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[3]),
    .en(al_1ce50ae3),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_ab2a7f1[3]));
  AL_DFF_X al_ad993ec1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[4]),
    .en(al_1ce50ae3),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_ab2a7f1[4]));
  AL_DFF_X al_2f6f2115 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[5]),
    .en(al_1ce50ae3),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_ab2a7f1[5]));
  AL_DFF_X al_11816c09 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[6]),
    .en(al_1ce50ae3),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_ab2a7f1[6]));
  AL_DFF_X al_dcbc3968 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[7]),
    .en(al_1ce50ae3),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_ab2a7f1[7]));
  AL_DFF_X al_5955dd2f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[8]),
    .en(al_1ce50ae3),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_ab2a7f1[8]));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff00f0f0ccccaaaa))
    al_55de7079 (
    .a(al_cd0aa0ee[0]),
    .b(al_25215c55[0]),
    .c(al_7808e039[0]),
    .d(al_a9406400),
    .e(al_82716c38[4]),
    .f(al_82716c38[5]),
    .o(al_f3899d20));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    al_1e122fd9 (
    .a(al_9b4eaefc[0]),
    .b(al_a0f12bef[0]),
    .c(al_868a1cad[0]),
    .d(al_82716c38[4]),
    .e(al_82716c38[5]),
    .o(al_1ca6a854));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfff30f5ffff3ff5f))
    al_d061d114 (
    .a(al_4096d0c7[0]),
    .b(al_ab2a7f1[0]),
    .c(al_82716c38[4]),
    .d(al_82716c38[5]),
    .e(al_82716c38[6]),
    .f(al_89a4ecab[0]),
    .o(al_d439eb63));
  AL_MAP_LUT6 #(
    .EQN("(D*~(~(~C*~(A)*~(E)+~C*A*~(E)+~(~C)*A*E+~C*A*E)*~(B)*~(F)+~(~C*~(A)*~(E)+~C*A*~(E)+~(~C)*A*E+~C*A*E)*B*~(F)+~(~(~C*~(A)*~(E)+~C*A*~(E)+~(~C)*A*E+~C*A*E))*B*F+~(~C*~(A)*~(E)+~C*A*~(E)+~(~C)*A*E+~C*A*E)*B*F))"),
    .INIT(64'h33003300aa000f00))
    al_18a51977 (
    .a(al_f3899d20),
    .b(al_d439eb63),
    .c(al_1ca6a854),
    .d(al_711bc49b),
    .e(al_82716c38[6]),
    .f(al_82716c38[7]),
    .o(al_492d1bb8[0]));
  AL_MAP_LUT6 #(
    .EQN("(~F*(A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E))"),
    .INIT(64'h00000000f0ccaa00))
    al_df9ca8e7 (
    .a(al_9b4eaefc[10]),
    .b(al_a0f12bef[10]),
    .c(al_868a1cad[10]),
    .d(al_82716c38[4]),
    .e(al_82716c38[5]),
    .f(al_82716c38[6]),
    .o(al_1e5502f4));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hfd3ffdff))
    al_b95b8ef3 (
    .a(al_ab2a7f1[10]),
    .b(al_82716c38[4]),
    .c(al_82716c38[5]),
    .d(al_82716c38[6]),
    .e(al_89a4ecab[10]),
    .o(al_2c28807a));
  AL_MAP_LUT6 #(
    .EQN("(C*~((~A*~(E*D))*~(B)*~(F)+(~A*~(E*D))*B*~(F)+~((~A*~(E*D)))*B*F+(~A*~(E*D))*B*F))"),
    .INIT(64'h30303030f0a0a0a0))
    al_7d38087d (
    .a(al_1e5502f4),
    .b(al_2c28807a),
    .c(al_711bc49b),
    .d(al_f751b948),
    .e(al_cd0aa0ee[10]),
    .f(al_82716c38[7]),
    .o(al_492d1bb8[10]));
  AL_MAP_LUT6 #(
    .EQN("(~F*(A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E))"),
    .INIT(64'h00000000f0ccaa00))
    al_8cb4e505 (
    .a(al_9b4eaefc[11]),
    .b(al_a0f12bef[11]),
    .c(al_868a1cad[11]),
    .d(al_82716c38[4]),
    .e(al_82716c38[5]),
    .f(al_82716c38[6]),
    .o(al_ccb46709));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hfd3ffdff))
    al_1b9c7863 (
    .a(al_ab2a7f1[11]),
    .b(al_82716c38[4]),
    .c(al_82716c38[5]),
    .d(al_82716c38[6]),
    .e(al_89a4ecab[11]),
    .o(al_f1c0edfa));
  AL_MAP_LUT6 #(
    .EQN("(C*~((~A*~(E*D))*~(B)*~(F)+(~A*~(E*D))*B*~(F)+~((~A*~(E*D)))*B*F+(~A*~(E*D))*B*F))"),
    .INIT(64'h30303030f0a0a0a0))
    al_a6a7777b (
    .a(al_ccb46709),
    .b(al_f1c0edfa),
    .c(al_711bc49b),
    .d(al_f751b948),
    .e(al_cd0aa0ee[11]),
    .f(al_82716c38[7]),
    .o(al_492d1bb8[11]));
  AL_MAP_LUT6 #(
    .EQN("(~F*(A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E))"),
    .INIT(64'h00000000f0ccaa00))
    al_7a83ee8e (
    .a(al_9b4eaefc[12]),
    .b(al_a0f12bef[12]),
    .c(al_868a1cad[12]),
    .d(al_82716c38[4]),
    .e(al_82716c38[5]),
    .f(al_82716c38[6]),
    .o(al_99b7d851));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hfd3ffdff))
    al_446a4d33 (
    .a(al_ab2a7f1[12]),
    .b(al_82716c38[4]),
    .c(al_82716c38[5]),
    .d(al_82716c38[6]),
    .e(al_89a4ecab[12]),
    .o(al_b945c2ed));
  AL_MAP_LUT6 #(
    .EQN("(C*~((~A*~(E*D))*~(B)*~(F)+(~A*~(E*D))*B*~(F)+~((~A*~(E*D)))*B*F+(~A*~(E*D))*B*F))"),
    .INIT(64'h30303030f0a0a0a0))
    al_196dabb6 (
    .a(al_99b7d851),
    .b(al_b945c2ed),
    .c(al_711bc49b),
    .d(al_f751b948),
    .e(al_cd0aa0ee[12]),
    .f(al_82716c38[7]),
    .o(al_492d1bb8[12]));
  AL_MAP_LUT6 #(
    .EQN("(~F*(A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E))"),
    .INIT(64'h00000000f0ccaa00))
    al_1968f3a2 (
    .a(al_9b4eaefc[13]),
    .b(al_a0f12bef[13]),
    .c(al_868a1cad[13]),
    .d(al_82716c38[4]),
    .e(al_82716c38[5]),
    .f(al_82716c38[6]),
    .o(al_337e2949));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hfd3ffdff))
    al_4184fc25 (
    .a(al_ab2a7f1[13]),
    .b(al_82716c38[4]),
    .c(al_82716c38[5]),
    .d(al_82716c38[6]),
    .e(al_89a4ecab[13]),
    .o(al_84914f7c));
  AL_MAP_LUT6 #(
    .EQN("(C*~((~A*~(E*D))*~(B)*~(F)+(~A*~(E*D))*B*~(F)+~((~A*~(E*D)))*B*F+(~A*~(E*D))*B*F))"),
    .INIT(64'h30303030f0a0a0a0))
    al_6804ce5d (
    .a(al_337e2949),
    .b(al_84914f7c),
    .c(al_711bc49b),
    .d(al_f751b948),
    .e(al_cd0aa0ee[13]),
    .f(al_82716c38[7]),
    .o(al_492d1bb8[13]));
  AL_MAP_LUT6 #(
    .EQN("(~F*(A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E))"),
    .INIT(64'h00000000f0ccaa00))
    al_799d3b47 (
    .a(al_9b4eaefc[14]),
    .b(al_a0f12bef[14]),
    .c(al_868a1cad[14]),
    .d(al_82716c38[4]),
    .e(al_82716c38[5]),
    .f(al_82716c38[6]),
    .o(al_ec6037b6));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hfd3ffdff))
    al_85c68a3c (
    .a(al_ab2a7f1[14]),
    .b(al_82716c38[4]),
    .c(al_82716c38[5]),
    .d(al_82716c38[6]),
    .e(al_89a4ecab[14]),
    .o(al_8e038ddf));
  AL_MAP_LUT6 #(
    .EQN("(C*~((~A*~(E*D))*~(B)*~(F)+(~A*~(E*D))*B*~(F)+~((~A*~(E*D)))*B*F+(~A*~(E*D))*B*F))"),
    .INIT(64'h30303030f0a0a0a0))
    al_721969d6 (
    .a(al_ec6037b6),
    .b(al_8e038ddf),
    .c(al_711bc49b),
    .d(al_f751b948),
    .e(al_cd0aa0ee[14]),
    .f(al_82716c38[7]),
    .o(al_492d1bb8[14]));
  AL_MAP_LUT6 #(
    .EQN("(~F*(A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E))"),
    .INIT(64'h00000000f0ccaa00))
    al_98168bc3 (
    .a(al_9b4eaefc[15]),
    .b(al_a0f12bef[15]),
    .c(al_868a1cad[15]),
    .d(al_82716c38[4]),
    .e(al_82716c38[5]),
    .f(al_82716c38[6]),
    .o(al_452179e4));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hfd3ffdff))
    al_ff1aa41f (
    .a(al_ab2a7f1[15]),
    .b(al_82716c38[4]),
    .c(al_82716c38[5]),
    .d(al_82716c38[6]),
    .e(al_89a4ecab[15]),
    .o(al_64bdbb03));
  AL_MAP_LUT6 #(
    .EQN("(C*~((~A*~(E*D))*~(B)*~(F)+(~A*~(E*D))*B*~(F)+~((~A*~(E*D)))*B*F+(~A*~(E*D))*B*F))"),
    .INIT(64'h30303030f0a0a0a0))
    al_d6864341 (
    .a(al_452179e4),
    .b(al_64bdbb03),
    .c(al_711bc49b),
    .d(al_f751b948),
    .e(al_cd0aa0ee[15]),
    .f(al_82716c38[7]),
    .o(al_492d1bb8[15]));
  AL_MAP_LUT6 #(
    .EQN("(A*(B*~(C)*~(D)*E*~(F)+B*C*~(D)*E*~(F)+B*~(C)*D*E*~(F)+B*C*D*E*~(F)+~(B)*C*~(D)*~(E)*F+B*C*~(D)*~(E)*F+~(B)*C*D*~(E)*F+B*C*D*~(E)*F+~(B)*~(C)*D*E*F+B*~(C)*D*E*F+~(B)*C*D*E*F+B*C*D*E*F))"),
    .INIT(64'haa00a0a088880000))
    al_17c94eec (
    .a(al_b256aea1),
    .b(al_9b4eaefc[16]),
    .c(al_a0f12bef[16]),
    .d(al_868a1cad[16]),
    .e(al_82716c38[4]),
    .f(al_82716c38[5]),
    .o(al_492d1bb8[16]));
  AL_MAP_LUT6 #(
    .EQN("(A*(B*~(C)*~(D)*E*~(F)+B*C*~(D)*E*~(F)+B*~(C)*D*E*~(F)+B*C*D*E*~(F)+~(B)*C*~(D)*~(E)*F+B*C*~(D)*~(E)*F+~(B)*C*D*~(E)*F+B*C*D*~(E)*F+~(B)*~(C)*D*E*F+B*~(C)*D*E*F+~(B)*C*D*E*F+B*C*D*E*F))"),
    .INIT(64'haa00a0a088880000))
    al_81b6e698 (
    .a(al_b256aea1),
    .b(al_9b4eaefc[17]),
    .c(al_a0f12bef[17]),
    .d(al_868a1cad[17]),
    .e(al_82716c38[4]),
    .f(al_82716c38[5]),
    .o(al_492d1bb8[17]));
  AL_MAP_LUT6 #(
    .EQN("(A*(B*~(C)*~(D)*E*~(F)+B*C*~(D)*E*~(F)+B*~(C)*D*E*~(F)+B*C*D*E*~(F)+~(B)*C*~(D)*~(E)*F+B*C*~(D)*~(E)*F+~(B)*C*D*~(E)*F+B*C*D*~(E)*F+~(B)*~(C)*D*E*F+B*~(C)*D*E*F+~(B)*C*D*E*F+B*C*D*E*F))"),
    .INIT(64'haa00a0a088880000))
    al_88e44d71 (
    .a(al_b256aea1),
    .b(al_9b4eaefc[18]),
    .c(al_a0f12bef[18]),
    .d(al_868a1cad[18]),
    .e(al_82716c38[4]),
    .f(al_82716c38[5]),
    .o(al_492d1bb8[18]));
  AL_MAP_LUT6 #(
    .EQN("(A*(B*~(C)*~(D)*E*~(F)+B*C*~(D)*E*~(F)+B*~(C)*D*E*~(F)+B*C*D*E*~(F)+~(B)*C*~(D)*~(E)*F+B*C*~(D)*~(E)*F+~(B)*C*D*~(E)*F+B*C*D*~(E)*F+~(B)*~(C)*D*E*F+B*~(C)*D*E*F+~(B)*C*D*E*F+B*C*D*E*F))"),
    .INIT(64'haa00a0a088880000))
    al_d325422d (
    .a(al_b256aea1),
    .b(al_9b4eaefc[19]),
    .c(al_a0f12bef[19]),
    .d(al_868a1cad[19]),
    .e(al_82716c38[4]),
    .f(al_82716c38[5]),
    .o(al_492d1bb8[19]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff0f3355))
    al_dd98aa40 (
    .a(al_cd0aa0ee[1]),
    .b(al_25215c55[1]),
    .c(al_7808e039[1]),
    .d(al_82716c38[4]),
    .e(al_82716c38[5]),
    .o(al_986ad8e6));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    al_5040d912 (
    .a(al_9b4eaefc[1]),
    .b(al_a0f12bef[1]),
    .c(al_868a1cad[1]),
    .d(al_82716c38[4]),
    .e(al_82716c38[5]),
    .o(al_d0cbf8c4));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfff30f5ffff3ff5f))
    al_efc6af1f (
    .a(al_4096d0c7[1]),
    .b(al_ab2a7f1[1]),
    .c(al_82716c38[4]),
    .d(al_82716c38[5]),
    .e(al_82716c38[6]),
    .f(al_89a4ecab[1]),
    .o(al_a4119c94));
  AL_MAP_LUT6 #(
    .EQN("(D*~((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(A)*~(F)+(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*~(F)+~((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*A*F+(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*F))"),
    .INIT(64'h5500550033000f00))
    al_dc318389 (
    .a(al_a4119c94),
    .b(al_986ad8e6),
    .c(al_d0cbf8c4),
    .d(al_711bc49b),
    .e(al_82716c38[6]),
    .f(al_82716c38[7]),
    .o(al_492d1bb8[1]));
  AL_MAP_LUT6 #(
    .EQN("(A*(B*~(C)*~(D)*E*~(F)+B*C*~(D)*E*~(F)+B*~(C)*D*E*~(F)+B*C*D*E*~(F)+~(B)*C*~(D)*~(E)*F+B*C*~(D)*~(E)*F+~(B)*C*D*~(E)*F+B*C*D*~(E)*F+~(B)*~(C)*D*E*F+B*~(C)*D*E*F+~(B)*C*D*E*F+B*C*D*E*F))"),
    .INIT(64'haa00a0a088880000))
    al_fbc1456b (
    .a(al_b256aea1),
    .b(al_9b4eaefc[20]),
    .c(al_a0f12bef[20]),
    .d(al_868a1cad[20]),
    .e(al_82716c38[4]),
    .f(al_82716c38[5]),
    .o(al_492d1bb8[20]));
  AL_MAP_LUT6 #(
    .EQN("(A*(B*~(C)*~(D)*E*~(F)+B*C*~(D)*E*~(F)+B*~(C)*D*E*~(F)+B*C*D*E*~(F)+~(B)*C*~(D)*~(E)*F+B*C*~(D)*~(E)*F+~(B)*C*D*~(E)*F+B*C*D*~(E)*F+~(B)*~(C)*D*E*F+B*~(C)*D*E*F+~(B)*C*D*E*F+B*C*D*E*F))"),
    .INIT(64'haa00a0a088880000))
    al_fb582983 (
    .a(al_b256aea1),
    .b(al_9b4eaefc[21]),
    .c(al_a0f12bef[21]),
    .d(al_868a1cad[21]),
    .e(al_82716c38[4]),
    .f(al_82716c38[5]),
    .o(al_492d1bb8[21]));
  AL_MAP_LUT6 #(
    .EQN("(A*(B*~(C)*~(D)*E*~(F)+B*C*~(D)*E*~(F)+B*~(C)*D*E*~(F)+B*C*D*E*~(F)+~(B)*C*~(D)*~(E)*F+B*C*~(D)*~(E)*F+~(B)*C*D*~(E)*F+B*C*D*~(E)*F+~(B)*~(C)*D*E*F+B*~(C)*D*E*F+~(B)*C*D*E*F+B*C*D*E*F))"),
    .INIT(64'haa00a0a088880000))
    al_be91e82b (
    .a(al_b256aea1),
    .b(al_9b4eaefc[22]),
    .c(al_a0f12bef[22]),
    .d(al_868a1cad[22]),
    .e(al_82716c38[4]),
    .f(al_82716c38[5]),
    .o(al_492d1bb8[22]));
  AL_MAP_LUT6 #(
    .EQN("(A*(B*~(C)*~(D)*E*~(F)+B*C*~(D)*E*~(F)+B*~(C)*D*E*~(F)+B*C*D*E*~(F)+~(B)*C*~(D)*~(E)*F+B*C*~(D)*~(E)*F+~(B)*C*D*~(E)*F+B*C*D*~(E)*F+~(B)*~(C)*D*E*F+B*~(C)*D*E*F+~(B)*C*D*E*F+B*C*D*E*F))"),
    .INIT(64'haa00a0a088880000))
    al_da14aaf3 (
    .a(al_b256aea1),
    .b(al_9b4eaefc[23]),
    .c(al_a0f12bef[23]),
    .d(al_868a1cad[23]),
    .e(al_82716c38[4]),
    .f(al_82716c38[5]),
    .o(al_492d1bb8[23]));
  AL_MAP_LUT6 #(
    .EQN("(A*(B*~(C)*~(D)*E*~(F)+B*C*~(D)*E*~(F)+B*~(C)*D*E*~(F)+B*C*D*E*~(F)+~(B)*C*~(D)*~(E)*F+B*C*~(D)*~(E)*F+~(B)*C*D*~(E)*F+B*C*D*~(E)*F+~(B)*~(C)*D*E*F+B*~(C)*D*E*F+~(B)*C*D*E*F+B*C*D*E*F))"),
    .INIT(64'haa00a0a088880000))
    al_56acfe28 (
    .a(al_b256aea1),
    .b(al_9b4eaefc[24]),
    .c(al_a0f12bef[24]),
    .d(al_868a1cad[24]),
    .e(al_82716c38[4]),
    .f(al_82716c38[5]),
    .o(al_492d1bb8[24]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_2244b1ea (
    .a(al_711bc49b),
    .b(al_82716c38[6]),
    .c(al_82716c38[7]),
    .o(al_b256aea1));
  AL_MAP_LUT6 #(
    .EQN("(A*(B*~(C)*~(D)*E*~(F)+B*C*~(D)*E*~(F)+B*~(C)*D*E*~(F)+B*C*D*E*~(F)+~(B)*C*~(D)*~(E)*F+B*C*~(D)*~(E)*F+~(B)*C*D*~(E)*F+B*C*D*~(E)*F+~(B)*~(C)*D*E*F+B*~(C)*D*E*F+~(B)*C*D*E*F+B*C*D*E*F))"),
    .INIT(64'haa00a0a088880000))
    al_5c1eedfd (
    .a(al_b256aea1),
    .b(al_9b4eaefc[25]),
    .c(al_a0f12bef[25]),
    .d(al_868a1cad[25]),
    .e(al_82716c38[4]),
    .f(al_82716c38[5]),
    .o(al_492d1bb8[25]));
  AL_MAP_LUT6 #(
    .EQN("(A*(B*~(C)*~(D)*E*~(F)+B*C*~(D)*E*~(F)+B*~(C)*D*E*~(F)+B*C*D*E*~(F)+~(B)*C*~(D)*~(E)*F+B*C*~(D)*~(E)*F+~(B)*C*D*~(E)*F+B*C*D*~(E)*F+~(B)*~(C)*D*E*F+B*~(C)*D*E*F+~(B)*C*D*E*F+B*C*D*E*F))"),
    .INIT(64'haa00a0a088880000))
    al_7cf92660 (
    .a(al_b256aea1),
    .b(al_9b4eaefc[26]),
    .c(al_a0f12bef[26]),
    .d(al_868a1cad[26]),
    .e(al_82716c38[4]),
    .f(al_82716c38[5]),
    .o(al_492d1bb8[26]));
  AL_MAP_LUT6 #(
    .EQN("(A*(B*~(C)*~(D)*E*~(F)+B*C*~(D)*E*~(F)+B*~(C)*D*E*~(F)+B*C*D*E*~(F)+~(B)*C*~(D)*~(E)*F+B*C*~(D)*~(E)*F+~(B)*C*D*~(E)*F+B*C*D*~(E)*F+~(B)*~(C)*D*E*F+B*~(C)*D*E*F+~(B)*C*D*E*F+B*C*D*E*F))"),
    .INIT(64'haa00a0a088880000))
    al_3bce26c2 (
    .a(al_b256aea1),
    .b(al_9b4eaefc[27]),
    .c(al_a0f12bef[27]),
    .d(al_868a1cad[27]),
    .e(al_82716c38[4]),
    .f(al_82716c38[5]),
    .o(al_492d1bb8[27]));
  AL_MAP_LUT6 #(
    .EQN("(A*(B*~(C)*~(D)*E*~(F)+B*C*~(D)*E*~(F)+B*~(C)*D*E*~(F)+B*C*D*E*~(F)+~(B)*C*~(D)*~(E)*F+B*C*~(D)*~(E)*F+~(B)*C*D*~(E)*F+B*C*D*~(E)*F+~(B)*~(C)*D*E*F+B*~(C)*D*E*F+~(B)*C*D*E*F+B*C*D*E*F))"),
    .INIT(64'haa00a0a088880000))
    al_e133b3a2 (
    .a(al_b256aea1),
    .b(al_9b4eaefc[28]),
    .c(al_a0f12bef[28]),
    .d(al_868a1cad[28]),
    .e(al_82716c38[4]),
    .f(al_82716c38[5]),
    .o(al_492d1bb8[28]));
  AL_MAP_LUT6 #(
    .EQN("(A*(B*~(C)*~(D)*E*~(F)+B*C*~(D)*E*~(F)+B*~(C)*D*E*~(F)+B*C*D*E*~(F)+~(B)*C*~(D)*~(E)*F+B*C*~(D)*~(E)*F+~(B)*C*D*~(E)*F+B*C*D*~(E)*F+~(B)*~(C)*D*E*F+B*~(C)*D*E*F+~(B)*C*D*E*F+B*C*D*E*F))"),
    .INIT(64'haa00a0a088880000))
    al_232bd57a (
    .a(al_b256aea1),
    .b(al_9b4eaefc[29]),
    .c(al_a0f12bef[29]),
    .d(al_868a1cad[29]),
    .e(al_82716c38[4]),
    .f(al_82716c38[5]),
    .o(al_492d1bb8[29]));
  AL_MAP_LUT6 #(
    .EQN("(~F*(A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E))"),
    .INIT(64'h00000000f0ccaa00))
    al_8ad561d5 (
    .a(al_9b4eaefc[2]),
    .b(al_a0f12bef[2]),
    .c(al_868a1cad[2]),
    .d(al_82716c38[4]),
    .e(al_82716c38[5]),
    .f(al_82716c38[6]),
    .o(al_19219cae));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfff30f5ffff3ff5f))
    al_e73ea44c (
    .a(al_4096d0c7[2]),
    .b(al_ab2a7f1[2]),
    .c(al_82716c38[4]),
    .d(al_82716c38[5]),
    .e(al_82716c38[6]),
    .f(al_89a4ecab[2]),
    .o(al_31650bb3));
  AL_MAP_LUT6 #(
    .EQN("(C*~((~A*~(E*D))*~(B)*~(F)+(~A*~(E*D))*B*~(F)+~((~A*~(E*D)))*B*F+(~A*~(E*D))*B*F))"),
    .INIT(64'h30303030f0a0a0a0))
    al_cc9357f4 (
    .a(al_19219cae),
    .b(al_31650bb3),
    .c(al_711bc49b),
    .d(al_f751b948),
    .e(al_cd0aa0ee[2]),
    .f(al_82716c38[7]),
    .o(al_492d1bb8[2]));
  AL_MAP_LUT6 #(
    .EQN("(A*(B*~(C)*~(D)*E*~(F)+B*C*~(D)*E*~(F)+B*~(C)*D*E*~(F)+B*C*D*E*~(F)+~(B)*C*~(D)*~(E)*F+B*C*~(D)*~(E)*F+~(B)*C*D*~(E)*F+B*C*D*~(E)*F+~(B)*~(C)*D*E*F+B*~(C)*D*E*F+~(B)*C*D*E*F+B*C*D*E*F))"),
    .INIT(64'haa00a0a088880000))
    al_1b32c3f8 (
    .a(al_b256aea1),
    .b(al_9b4eaefc[30]),
    .c(al_a0f12bef[30]),
    .d(al_868a1cad[30]),
    .e(al_82716c38[4]),
    .f(al_82716c38[5]),
    .o(al_492d1bb8[30]));
  AL_MAP_LUT6 #(
    .EQN("(A*(B*~(C)*~(D)*E*~(F)+B*C*~(D)*E*~(F)+B*~(C)*D*E*~(F)+B*C*D*E*~(F)+~(B)*C*~(D)*~(E)*F+B*C*~(D)*~(E)*F+~(B)*C*D*~(E)*F+B*C*D*~(E)*F+~(B)*~(C)*D*E*F+B*~(C)*D*E*F+~(B)*C*D*E*F+B*C*D*E*F))"),
    .INIT(64'haa00a0a088880000))
    al_61470d6e (
    .a(al_b256aea1),
    .b(al_9b4eaefc[31]),
    .c(al_a0f12bef[31]),
    .d(al_868a1cad[31]),
    .e(al_82716c38[4]),
    .f(al_82716c38[5]),
    .o(al_492d1bb8[31]));
  AL_MAP_LUT6 #(
    .EQN("(~F*(A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E))"),
    .INIT(64'h00000000f0ccaa00))
    al_2e10fd26 (
    .a(al_9b4eaefc[3]),
    .b(al_a0f12bef[3]),
    .c(al_868a1cad[3]),
    .d(al_82716c38[4]),
    .e(al_82716c38[5]),
    .f(al_82716c38[6]),
    .o(al_97f75483));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfff30f5ffff3ff5f))
    al_2b136760 (
    .a(al_4096d0c7[3]),
    .b(al_ab2a7f1[3]),
    .c(al_82716c38[4]),
    .d(al_82716c38[5]),
    .e(al_82716c38[6]),
    .f(al_89a4ecab[3]),
    .o(al_df62d485));
  AL_MAP_LUT6 #(
    .EQN("(C*~((~A*~(E*D))*~(B)*~(F)+(~A*~(E*D))*B*~(F)+~((~A*~(E*D)))*B*F+(~A*~(E*D))*B*F))"),
    .INIT(64'h30303030f0a0a0a0))
    al_b109267b (
    .a(al_97f75483),
    .b(al_df62d485),
    .c(al_711bc49b),
    .d(al_f751b948),
    .e(al_cd0aa0ee[3]),
    .f(al_82716c38[7]),
    .o(al_492d1bb8[3]));
  AL_MAP_LUT6 #(
    .EQN("(~F*(A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E))"),
    .INIT(64'h00000000f0ccaa00))
    al_db80aa6c (
    .a(al_9b4eaefc[4]),
    .b(al_a0f12bef[4]),
    .c(al_868a1cad[4]),
    .d(al_82716c38[4]),
    .e(al_82716c38[5]),
    .f(al_82716c38[6]),
    .o(al_1a3cae1d));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfff30f5ffff3ff5f))
    al_63d71e59 (
    .a(al_4096d0c7[4]),
    .b(al_ab2a7f1[4]),
    .c(al_82716c38[4]),
    .d(al_82716c38[5]),
    .e(al_82716c38[6]),
    .f(al_89a4ecab[4]),
    .o(al_60cada77));
  AL_MAP_LUT6 #(
    .EQN("(C*~((~A*~(E*D))*~(B)*~(F)+(~A*~(E*D))*B*~(F)+~((~A*~(E*D)))*B*F+(~A*~(E*D))*B*F))"),
    .INIT(64'h30303030f0a0a0a0))
    al_298047a1 (
    .a(al_1a3cae1d),
    .b(al_60cada77),
    .c(al_711bc49b),
    .d(al_f751b948),
    .e(al_cd0aa0ee[4]),
    .f(al_82716c38[7]),
    .o(al_492d1bb8[4]));
  AL_MAP_LUT6 #(
    .EQN("(~F*(A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E))"),
    .INIT(64'h00000000f0ccaa00))
    al_4aadee06 (
    .a(al_9b4eaefc[5]),
    .b(al_a0f12bef[5]),
    .c(al_868a1cad[5]),
    .d(al_82716c38[4]),
    .e(al_82716c38[5]),
    .f(al_82716c38[6]),
    .o(al_f817c39d));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfff30f5ffff3ff5f))
    al_a9123b67 (
    .a(al_4096d0c7[5]),
    .b(al_ab2a7f1[5]),
    .c(al_82716c38[4]),
    .d(al_82716c38[5]),
    .e(al_82716c38[6]),
    .f(al_89a4ecab[5]),
    .o(al_1041edd0));
  AL_MAP_LUT6 #(
    .EQN("(C*~((~A*~(E*D))*~(B)*~(F)+(~A*~(E*D))*B*~(F)+~((~A*~(E*D)))*B*F+(~A*~(E*D))*B*F))"),
    .INIT(64'h30303030f0a0a0a0))
    al_e5330f41 (
    .a(al_f817c39d),
    .b(al_1041edd0),
    .c(al_711bc49b),
    .d(al_f751b948),
    .e(al_cd0aa0ee[5]),
    .f(al_82716c38[7]),
    .o(al_492d1bb8[5]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_167760d4 (
    .a(al_82716c38[0]),
    .b(al_82716c38[1]),
    .c(al_82716c38[2]),
    .d(al_82716c38[3]),
    .o(al_711bc49b));
  AL_MAP_LUT6 #(
    .EQN("(C*~((~B*~(E*D))*~(A)*~(F)+(~B*~(E*D))*A*~(F)+~((~B*~(E*D)))*A*F+(~B*~(E*D))*A*F))"),
    .INIT(64'h50505050f0c0c0c0))
    al_b270e2ba (
    .a(al_7e094735),
    .b(al_36697857),
    .c(al_711bc49b),
    .d(al_f751b948),
    .e(al_cd0aa0ee[6]),
    .f(al_82716c38[7]),
    .o(al_492d1bb8[6]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_9ec140ec (
    .a(al_82716c38[4]),
    .b(al_82716c38[5]),
    .c(al_82716c38[6]),
    .o(al_f751b948));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_62071db2 (
    .a(al_4096d0c7[0]),
    .b(al_4096d0c7[1]),
    .c(al_4096d0c7[2]),
    .d(al_4096d0c7[3]),
    .e(al_4096d0c7[4]),
    .f(al_4096d0c7[5]),
    .o(al_37d9882e));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_30e3aa9c (
    .a(al_37d9882e),
    .b(al_4096d0c7[6]),
    .o(al_fd9c8287));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfff30f5ffff3ff5f))
    al_853ba5e9 (
    .a(al_fd9c8287),
    .b(al_ab2a7f1[6]),
    .c(al_82716c38[4]),
    .d(al_82716c38[5]),
    .e(al_82716c38[6]),
    .f(al_89a4ecab[6]),
    .o(al_7e094735));
  AL_MAP_LUT6 #(
    .EQN("(~F*(A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E))"),
    .INIT(64'h00000000f0ccaa00))
    al_df0f2b37 (
    .a(al_9b4eaefc[6]),
    .b(al_a0f12bef[6]),
    .c(al_868a1cad[6]),
    .d(al_82716c38[4]),
    .e(al_82716c38[5]),
    .f(al_82716c38[6]),
    .o(al_36697857));
  AL_MAP_LUT6 #(
    .EQN("(~F*(A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E))"),
    .INIT(64'h00000000f0ccaa00))
    al_cbeea0a0 (
    .a(al_9b4eaefc[7]),
    .b(al_a0f12bef[7]),
    .c(al_868a1cad[7]),
    .d(al_82716c38[4]),
    .e(al_82716c38[5]),
    .f(al_82716c38[6]),
    .o(al_9e512d7f));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hfd3ffdff))
    al_f0f0cfb9 (
    .a(al_ab2a7f1[7]),
    .b(al_82716c38[4]),
    .c(al_82716c38[5]),
    .d(al_82716c38[6]),
    .e(al_89a4ecab[7]),
    .o(al_d889aa1d));
  AL_MAP_LUT6 #(
    .EQN("(C*~((~A*~(E*D))*~(B)*~(F)+(~A*~(E*D))*B*~(F)+~((~A*~(E*D)))*B*F+(~A*~(E*D))*B*F))"),
    .INIT(64'h30303030f0a0a0a0))
    al_b88e8ebd (
    .a(al_9e512d7f),
    .b(al_d889aa1d),
    .c(al_711bc49b),
    .d(al_f751b948),
    .e(al_cd0aa0ee[7]),
    .f(al_82716c38[7]),
    .o(al_492d1bb8[7]));
  AL_MAP_LUT6 #(
    .EQN("(~F*(A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E))"),
    .INIT(64'h00000000f0ccaa00))
    al_db7855fc (
    .a(al_9b4eaefc[8]),
    .b(al_a0f12bef[8]),
    .c(al_868a1cad[8]),
    .d(al_82716c38[4]),
    .e(al_82716c38[5]),
    .f(al_82716c38[6]),
    .o(al_45b5d05e));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hfd3ffdff))
    al_b7a8370b (
    .a(al_ab2a7f1[8]),
    .b(al_82716c38[4]),
    .c(al_82716c38[5]),
    .d(al_82716c38[6]),
    .e(al_89a4ecab[8]),
    .o(al_9f0f27fb));
  AL_MAP_LUT6 #(
    .EQN("(C*~((~A*~(E*D))*~(B)*~(F)+(~A*~(E*D))*B*~(F)+~((~A*~(E*D)))*B*F+(~A*~(E*D))*B*F))"),
    .INIT(64'h30303030f0a0a0a0))
    al_beeb510 (
    .a(al_45b5d05e),
    .b(al_9f0f27fb),
    .c(al_711bc49b),
    .d(al_f751b948),
    .e(al_cd0aa0ee[8]),
    .f(al_82716c38[7]),
    .o(al_492d1bb8[8]));
  AL_MAP_LUT6 #(
    .EQN("(~F*(A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E))"),
    .INIT(64'h00000000f0ccaa00))
    al_32b67c5f (
    .a(al_9b4eaefc[9]),
    .b(al_a0f12bef[9]),
    .c(al_868a1cad[9]),
    .d(al_82716c38[4]),
    .e(al_82716c38[5]),
    .f(al_82716c38[6]),
    .o(al_153ccbd8));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hfd3ffdff))
    al_d078e817 (
    .a(al_ab2a7f1[9]),
    .b(al_82716c38[4]),
    .c(al_82716c38[5]),
    .d(al_82716c38[6]),
    .e(al_89a4ecab[9]),
    .o(al_eae41b9d));
  AL_MAP_LUT6 #(
    .EQN("(C*~((~A*~(E*D))*~(B)*~(F)+(~A*~(E*D))*B*~(F)+~((~A*~(E*D)))*B*F+(~A*~(E*D))*B*F))"),
    .INIT(64'h30303030f0a0a0a0))
    al_7b8b16c9 (
    .a(al_153ccbd8),
    .b(al_eae41b9d),
    .c(al_711bc49b),
    .d(al_f751b948),
    .e(al_cd0aa0ee[9]),
    .f(al_82716c38[7]),
    .o(al_492d1bb8[9]));
  AL_DFF_X al_9aa6335b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_d016a646),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7968b2a5));
  AL_MAP_LUT6 #(
    .EQN("(~B*(D*~(A)*~((F*E*~C))+D*A*~((F*E*~C))+~(D)*A*(F*E*~C)+D*A*(F*E*~C)))"),
    .INIT(64'h3202330033003300))
    al_1a0e74b0 (
    .a(al_fd9c8287),
    .b(al_81344cef),
    .c(al_6b181c0),
    .d(al_7968b2a5),
    .e(al_c9bfee53),
    .f(al_7c711acd),
    .o(al_d016a646));
  AL_DFF_X al_28356984 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_6b181c0),
    .en(1'b1),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_7c711acd));
  AL_DFF_X al_4cfc1aa4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(mdio_in),
    .en(1'b1),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_14e5d384));
  AL_DFF_X al_5940691 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_14e5d384),
    .en(1'b1),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_c6d1dc18));
  AL_DFF_X al_682a90fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9befeaf3),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mdio_out));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+A*~(B)*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'haaaaccccf0f0ff00))
    al_ac1a8ed9 (
    .a(al_523025ae[4]),
    .b(al_523025ae[5]),
    .c(al_523025ae[6]),
    .d(al_523025ae[7]),
    .e(al_ec1f16c4[0]),
    .f(al_ec1f16c4[1]),
    .o(al_62e089bb));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+A*~(B)*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hf0f0aaaacccc00ff))
    al_478cd5f5 (
    .a(al_33409841),
    .b(al_62e089bb),
    .c(al_eb828cf9),
    .d(al_6dd1a6b),
    .e(al_ec1f16c4[2]),
    .f(al_ec1f16c4[3]),
    .o(al_4db525a4));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+A*~(B)*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'haaaaccccf0f0ff00))
    al_a0feafdb (
    .a(al_ab2a7f1[8]),
    .b(al_ab2a7f1[9]),
    .c(al_ab2a7f1[10]),
    .d(al_ab2a7f1[11]),
    .e(al_ec1f16c4[0]),
    .f(al_ec1f16c4[1]),
    .o(al_75328a30));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+A*~(B)*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'haaaaccccf0f0ff00))
    al_74d68817 (
    .a(al_ab2a7f1[0]),
    .b(al_ab2a7f1[1]),
    .c(al_ab2a7f1[2]),
    .d(al_ab2a7f1[3]),
    .e(al_ec1f16c4[0]),
    .f(al_ec1f16c4[1]),
    .o(al_47962165));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+A*~(B)*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'haaaaccccf0f0ff00))
    al_14550e7f (
    .a(al_ab2a7f1[12]),
    .b(al_ab2a7f1[13]),
    .c(al_ab2a7f1[14]),
    .d(al_ab2a7f1[15]),
    .e(al_ec1f16c4[0]),
    .f(al_ec1f16c4[1]),
    .o(al_53937ca8));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+A*~(B)*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+A*~(B)*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+A*B*~(C)*D*E*F+A*~(B)*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'haaaaccccf0f0ff00))
    al_1702f10a (
    .a(al_ab2a7f1[4]),
    .b(al_ab2a7f1[5]),
    .c(al_ab2a7f1[6]),
    .d(al_ab2a7f1[7]),
    .e(al_ec1f16c4[0]),
    .f(al_ec1f16c4[1]),
    .o(al_6bda5d58));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+A*~(B)*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hccccff00aaaaf0f0))
    al_31d78843 (
    .a(al_75328a30),
    .b(al_47962165),
    .c(al_53937ca8),
    .d(al_6bda5d58),
    .e(al_ec1f16c4[2]),
    .f(al_ec1f16c4[3]),
    .o(al_c3f8fcfd));
  AL_MAP_LUT4 #(
    .EQN("(D*~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h5300))
    al_260dc47e (
    .a(al_c3f8fcfd),
    .b(al_4db525a4),
    .c(al_ec1f16c4[4]),
    .d(al_ec1f16c4[5]),
    .o(al_ca75b795));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(~D*~(A)*~((E*~C))+~D*A*~((E*~C))+~(~D)*A*(E*~C)+~D*A*(E*~C)))"),
    .INIT(32'h31013300))
    al_af973ba5 (
    .a(al_ca75b795),
    .b(al_81344cef),
    .c(al_6b181c0),
    .d(mdio_out),
    .e(al_7c711acd),
    .o(al_9befeaf3));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hccccf0f0ff00aaaa))
    al_7aa5978 (
    .a(al_523025ae[3]),
    .b(al_523025ae[10]),
    .c(al_523025ae[11]),
    .d(al_523025ae[12]),
    .e(al_ec1f16c4[0]),
    .f(al_ec1f16c4[1]),
    .o(al_33409841));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    al_43c93f9 (
    .a(al_523025ae[8]),
    .b(al_523025ae[9]),
    .c(al_ec1f16c4[0]),
    .d(al_ec1f16c4[1]),
    .o(al_eb828cf9));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h530f))
    al_27cfd3eb (
    .a(al_523025ae[1]),
    .b(al_523025ae[2]),
    .c(al_ec1f16c4[0]),
    .d(al_ec1f16c4[1]),
    .o(al_6dd1a6b));
  AL_DFF_X al_e07284fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_d376e8f0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mdio_oen));
  AL_MAP_LUT6 #(
    .EQN("(F*A*~(~E*~(D*C*B)))"),
    .INIT(64'haaaa800000000000))
    al_fdbf8295 (
    .a(al_523025ae[2]),
    .b(al_ec1f16c4[1]),
    .c(al_ec1f16c4[2]),
    .d(al_ec1f16c4[3]),
    .e(al_ec1f16c4[4]),
    .f(al_ec1f16c4[5]),
    .o(al_e25f50ab));
  AL_MAP_LUT6 #(
    .EQN("~(~B*(~D*~((~E*~A))*~((F*~C))+~D*(~E*~A)*~((F*~C))+~(~D)*(~E*~A)*(F*~C)+~D*(~E*~A)*(F*~C)))"),
    .INIT(64'hffcffeceffccffcc))
    al_43746dcb (
    .a(al_e25f50ab),
    .b(al_81344cef),
    .c(al_6b181c0),
    .d(mdio_oen),
    .e(al_c9bfee53),
    .f(al_7c711acd),
    .o(al_d376e8f0));
  AL_DFF_X al_56f2a50b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_2dc26b59),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c9bfee53));
  AL_MAP_LUT6 #(
    .EQN("~(~C*(~(A)*~(B)*~((E*D))*~(F)+A*~(B)*~((E*D))*~(F)+~(A)*B*~((E*D))*~(F)+~(A)*~(B)*(E*D)*~(F)+A*~(B)*(E*D)*~(F)+~(A)*B*(E*D)*~(F)+~(A)*B*(E*D)*F))"),
    .INIT(64'hfbfffffff8f8f8f8))
    al_dc8a8e0a (
    .a(al_6a1aebd1),
    .b(al_3cbc9279),
    .c(al_81344cef),
    .d(al_8587a543),
    .e(al_7968b2a5),
    .f(al_c9bfee53),
    .o(al_2dc26b59));
  AL_DFF_X al_f96bcb86 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_314de0e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec1f16c4[0]));
  AL_DFF_X al_d7c373fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_84d6d5e6),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec1f16c4[1]));
  AL_DFF_X al_b9c823d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_70a55548),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec1f16c4[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_247db07f (
    .a(al_ec1f16c4[0]),
    .b(al_ec1f16c4[1]),
    .c(al_ec1f16c4[2]),
    .o(al_a511ca2d));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_f940d705 (
    .a(al_a511ca2d),
    .b(al_ec1f16c4[3]),
    .c(al_ec1f16c4[4]),
    .o(al_60c51ee3));
  AL_DFF_X al_e6c73aa1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_a51b1b3a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec1f16c4[3]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_a45bddfb (
    .a(al_6b181c0),
    .b(al_7c711acd),
    .o(al_3cbc9279));
  AL_MAP_LUT5 #(
    .EQN("(~B*(A*~(C)*D*~(E)+~(A)*~(C)*~(D)*E+A*~(C)*~(D)*E+~(A)*C*~(D)*E+~(A)*~(C)*D*E+~(A)*C*D*E))"),
    .INIT(32'h11130200))
    al_eab90def (
    .a(al_3cbc9279),
    .b(al_81344cef),
    .c(al_c9bfee53),
    .d(al_ec1f16c4[0]),
    .e(al_ec1f16c4[1]),
    .o(al_84d6d5e6));
  AL_MAP_LUT4 #(
    .EQN("(~B*(A*~(C)*~(D)+~(A)*~(C)*D+~(A)*C*D))"),
    .INIT(16'h1102))
    al_f2b86327 (
    .a(al_3cbc9279),
    .b(al_81344cef),
    .c(al_c9bfee53),
    .d(al_ec1f16c4[0]),
    .o(al_314de0e));
  AL_MAP_LUT6 #(
    .EQN("(~B*(A*~(C)*(E*D)*~(F)+~(A)*~(C)*~((E*D))*F+A*~(C)*~((E*D))*F+~(A)*C*~((E*D))*F+~(A)*~(C)*(E*D)*F+~(A)*C*(E*D)*F))"),
    .INIT(64'h1113131302000000))
    al_803f894 (
    .a(al_3cbc9279),
    .b(al_81344cef),
    .c(al_c9bfee53),
    .d(al_ec1f16c4[0]),
    .e(al_ec1f16c4[1]),
    .f(al_ec1f16c4[2]),
    .o(al_70a55548));
  AL_MAP_LUT5 #(
    .EQN("(~C*(A*B*~(D)*~(E)+~(A)*~(B)*~(D)*E+A*~(B)*~(D)*E+~(A)*B*~(D)*E+~(A)*~(B)*D*E+A*~(B)*D*E))"),
    .INIT(32'h03070008))
    al_c21842e7 (
    .a(al_a511ca2d),
    .b(al_3cbc9279),
    .c(al_81344cef),
    .d(al_c9bfee53),
    .e(al_ec1f16c4[3]),
    .o(al_a51b1b3a));
  AL_MAP_LUT6 #(
    .EQN("(~C*(B*~(D)*(E*A)*~(F)+~(B)*~(D)*~((E*A))*F+B*~(D)*~((E*A))*F+~(B)*D*~((E*A))*F+~(B)*~(D)*(E*A)*F+~(B)*D*(E*A)*F))"),
    .INIT(64'h0307030f00080000))
    al_39cbfd77 (
    .a(al_a511ca2d),
    .b(al_3cbc9279),
    .c(al_81344cef),
    .d(al_c9bfee53),
    .e(al_ec1f16c4[3]),
    .f(al_ec1f16c4[4]),
    .o(al_acb683b9));
  AL_MAP_LUT5 #(
    .EQN("(~C*(A*B*~(D)*~(E)+~(A)*~(B)*~(D)*E+A*~(B)*~(D)*E+~(A)*B*~(D)*E+~(A)*~(B)*D*E+A*~(B)*D*E))"),
    .INIT(32'h03070008))
    al_985e3639 (
    .a(al_60c51ee3),
    .b(al_3cbc9279),
    .c(al_81344cef),
    .d(al_c9bfee53),
    .e(al_ec1f16c4[5]),
    .o(al_7f071305));
  AL_DFF_X al_41623954 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_acb683b9),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec1f16c4[4]));
  AL_DFF_X al_bc43eae0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_7f071305),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ec1f16c4[5]));
  AL_DFF_X al_c314d5c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_c53dc261),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_89a4ecab[0]));
  AL_DFF_X al_b09b0d1f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_2014d3d9),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_89a4ecab[9]));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F*~(C)*~((~E*D*A))+F*C*~((~E*D*A))+~(F)*C*(~E*D*A)+F*C*(~E*D*A)))"),
    .INIT(64'h3333313300002000))
    al_7466861d (
    .a(al_572dc31a),
    .b(al_81344cef),
    .c(al_c6d1dc18),
    .d(al_ec1f16c4[0]),
    .e(al_ec1f16c4[1]),
    .f(al_89a4ecab[14]),
    .o(al_48bec3d3));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F*~(C)*~((E*~D*A))+F*C*~((E*~D*A))+~(F)*C*(E*~D*A)+F*C*(E*~D*A)))"),
    .INIT(64'h3331333300200000))
    al_3d4d8dee (
    .a(al_572dc31a),
    .b(al_81344cef),
    .c(al_c6d1dc18),
    .d(al_ec1f16c4[0]),
    .e(al_ec1f16c4[1]),
    .f(al_89a4ecab[13]),
    .o(al_c1b912e));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F*~(C)*~((E*D*A))+F*C*~((E*D*A))+~(F)*C*(E*D*A)+F*C*(E*D*A)))"),
    .INIT(64'h3133333320000000))
    al_50a1f9f0 (
    .a(al_572dc31a),
    .b(al_81344cef),
    .c(al_c6d1dc18),
    .d(al_ec1f16c4[0]),
    .e(al_ec1f16c4[1]),
    .f(al_89a4ecab[12]),
    .o(al_aacd2311));
  AL_MAP_LUT5 #(
    .EQN("(~C*(E*~(D)*~((B*A))+E*D*~((B*A))+~(E)*D*(B*A)+E*D*(B*A)))"),
    .INIT(32'h0f070800))
    al_59caa487 (
    .a(al_6a1aebd1),
    .b(al_3cbc9279),
    .c(al_81344cef),
    .d(al_c6d1dc18),
    .e(al_89a4ecab[0]),
    .o(al_c53dc261));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    al_5b93e20f (
    .a(al_3cbc9279),
    .b(al_ec1f16c4[2]),
    .c(al_ec1f16c4[3]),
    .d(al_ec1f16c4[4]),
    .e(al_ec1f16c4[5]),
    .o(al_3b935332));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F*~(C)*~((E*~D*A))+F*C*~((E*~D*A))+~(F)*C*(E*~D*A)+F*C*(E*~D*A)))"),
    .INIT(64'h3331333300200000))
    al_44c533db (
    .a(al_3b935332),
    .b(al_81344cef),
    .c(al_c6d1dc18),
    .d(al_ec1f16c4[0]),
    .e(al_ec1f16c4[1]),
    .f(al_89a4ecab[1]),
    .o(al_e7834cb3));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F*~(C)*~((~E*D*A))+F*C*~((~E*D*A))+~(F)*C*(~E*D*A)+F*C*(~E*D*A)))"),
    .INIT(64'h3333313300002000))
    al_bf2b75a9 (
    .a(al_3b935332),
    .b(al_81344cef),
    .c(al_c6d1dc18),
    .d(al_ec1f16c4[0]),
    .e(al_ec1f16c4[1]),
    .f(al_89a4ecab[2]),
    .o(al_144281a5));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F*~(C)*~((~E*~D*A))+F*C*~((~E*~D*A))+~(F)*C*(~E*~D*A)+F*C*(~E*~D*A)))"),
    .INIT(64'h3333333100000020))
    al_32882e67 (
    .a(al_3b935332),
    .b(al_81344cef),
    .c(al_c6d1dc18),
    .d(al_ec1f16c4[0]),
    .e(al_ec1f16c4[1]),
    .f(al_89a4ecab[3]),
    .o(al_dcaf20fc));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*~B*A)"),
    .INIT(32'h20000000))
    al_ea21bc35 (
    .a(al_3cbc9279),
    .b(al_ec1f16c4[2]),
    .c(al_ec1f16c4[3]),
    .d(al_ec1f16c4[4]),
    .e(al_ec1f16c4[5]),
    .o(al_c68dfd58));
  AL_DFF_X al_4d8a64b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_39855db7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_89a4ecab[10]));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F*~(C)*~((E*D*A))+F*C*~((E*D*A))+~(F)*C*(E*D*A)+F*C*(E*D*A)))"),
    .INIT(64'h3133333320000000))
    al_b1cca85c (
    .a(al_c68dfd58),
    .b(al_81344cef),
    .c(al_c6d1dc18),
    .d(al_ec1f16c4[0]),
    .e(al_ec1f16c4[1]),
    .f(al_89a4ecab[4]),
    .o(al_ad53d9d0));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F*~(C)*~((E*~D*A))+F*C*~((E*~D*A))+~(F)*C*(E*~D*A)+F*C*(E*~D*A)))"),
    .INIT(64'h3331333300200000))
    al_95af5ed8 (
    .a(al_c68dfd58),
    .b(al_81344cef),
    .c(al_c6d1dc18),
    .d(al_ec1f16c4[0]),
    .e(al_ec1f16c4[1]),
    .f(al_89a4ecab[5]),
    .o(al_ffec892d));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F*~(C)*~((~E*D*A))+F*C*~((~E*D*A))+~(F)*C*(~E*D*A)+F*C*(~E*D*A)))"),
    .INIT(64'h3333313300002000))
    al_67296513 (
    .a(al_c68dfd58),
    .b(al_81344cef),
    .c(al_c6d1dc18),
    .d(al_ec1f16c4[0]),
    .e(al_ec1f16c4[1]),
    .f(al_89a4ecab[6]),
    .o(al_d24d858b));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F*~(C)*~((~E*~D*A))+F*C*~((~E*~D*A))+~(F)*C*(~E*~D*A)+F*C*(~E*~D*A)))"),
    .INIT(64'h3333333100000020))
    al_53f17a9b (
    .a(al_c68dfd58),
    .b(al_81344cef),
    .c(al_c6d1dc18),
    .d(al_ec1f16c4[0]),
    .e(al_ec1f16c4[1]),
    .f(al_89a4ecab[7]),
    .o(al_6400d4de));
  AL_MAP_LUT5 #(
    .EQN("(E*D*~C*B*A)"),
    .INIT(32'h08000000))
    al_cc9383ca (
    .a(al_3cbc9279),
    .b(al_ec1f16c4[2]),
    .c(al_ec1f16c4[3]),
    .d(al_ec1f16c4[4]),
    .e(al_ec1f16c4[5]),
    .o(al_4e8c0a64));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F*~(C)*~((E*D*A))+F*C*~((E*D*A))+~(F)*C*(E*D*A)+F*C*(E*D*A)))"),
    .INIT(64'h3133333320000000))
    al_b326f9b2 (
    .a(al_4e8c0a64),
    .b(al_81344cef),
    .c(al_c6d1dc18),
    .d(al_ec1f16c4[0]),
    .e(al_ec1f16c4[1]),
    .f(al_89a4ecab[8]),
    .o(al_e8e15f03));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F*~(C)*~((E*~D*A))+F*C*~((E*~D*A))+~(F)*C*(E*~D*A)+F*C*(E*~D*A)))"),
    .INIT(64'h3331333300200000))
    al_edc595ec (
    .a(al_4e8c0a64),
    .b(al_81344cef),
    .c(al_c6d1dc18),
    .d(al_ec1f16c4[0]),
    .e(al_ec1f16c4[1]),
    .f(al_89a4ecab[9]),
    .o(al_2014d3d9));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F*~(C)*~((~E*D*A))+F*C*~((~E*D*A))+~(F)*C*(~E*D*A)+F*C*(~E*D*A)))"),
    .INIT(64'h3333313300002000))
    al_b1cfecd (
    .a(al_4e8c0a64),
    .b(al_81344cef),
    .c(al_c6d1dc18),
    .d(al_ec1f16c4[0]),
    .e(al_ec1f16c4[1]),
    .f(al_89a4ecab[10]),
    .o(al_39855db7));
  AL_DFF_X al_7d1cc482 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_6230936a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_89a4ecab[11]));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F*~(C)*~((~E*~D*A))+F*C*~((~E*~D*A))+~(F)*C*(~E*~D*A)+F*C*(~E*~D*A)))"),
    .INIT(64'h3333333100000020))
    al_322c78ed (
    .a(al_4e8c0a64),
    .b(al_81344cef),
    .c(al_c6d1dc18),
    .d(al_ec1f16c4[0]),
    .e(al_ec1f16c4[1]),
    .f(al_89a4ecab[11]),
    .o(al_6230936a));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F*~(C)*~((~E*~D*A))+F*C*~((~E*~D*A))+~(F)*C*(~E*~D*A)+F*C*(~E*~D*A)))"),
    .INIT(64'h3333333100000020))
    al_62a975ef (
    .a(al_572dc31a),
    .b(al_81344cef),
    .c(al_c6d1dc18),
    .d(al_ec1f16c4[0]),
    .e(al_ec1f16c4[1]),
    .f(al_89a4ecab[15]),
    .o(al_751a5b13));
  AL_DFF_X al_3e2a87d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_aacd2311),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_89a4ecab[12]));
  AL_DFF_X al_177962f3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_c1b912e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_89a4ecab[13]));
  AL_DFF_X al_f33caacf (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_48bec3d3),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_89a4ecab[14]));
  AL_DFF_X al_e2030f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_751a5b13),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_89a4ecab[15]));
  AL_DFF_X al_f22402a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_e7834cb3),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_89a4ecab[1]));
  AL_DFF_X al_6014c805 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_144281a5),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_89a4ecab[2]));
  AL_DFF_X al_643d23fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_dcaf20fc),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_89a4ecab[3]));
  AL_DFF_X al_398e6346 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ad53d9d0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_89a4ecab[4]));
  AL_DFF_X al_bb42c111 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_ffec892d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_89a4ecab[5]));
  AL_DFF_X al_b769f9e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_d24d858b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_89a4ecab[6]));
  AL_DFF_X al_e0ca9824 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_6400d4de),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_89a4ecab[7]));
  AL_DFF_X al_2aa3963 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_e8e15f03),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_89a4ecab[8]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_36a6b003 (
    .a(al_60c51ee3),
    .b(al_ec1f16c4[5]),
    .o(al_6a1aebd1));
  AL_MAP_LUT5 #(
    .EQN("(E*D*~C*~B*A)"),
    .INIT(32'h02000000))
    al_6950fe3f (
    .a(al_3cbc9279),
    .b(al_ec1f16c4[2]),
    .c(al_ec1f16c4[3]),
    .d(al_ec1f16c4[4]),
    .e(al_ec1f16c4[5]),
    .o(al_572dc31a));
  AL_DFF_X al_21a36285 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_6a1aebd1),
    .en(1'b1),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_2b48f483));
  AL_DFF_X al_c28b1c09 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_2b48f483),
    .en(1'b1),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_841146bf));
  AL_DFF_X al_71730d86 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_af3abf3a),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_5772dfd3));
  AL_DFF_X al_8a745304 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_3e7ed8af),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_e2b7a540));
  AL_DFF_X al_37eb0453 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_cb74bfe8),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c5bc3747));
  AL_MAP_LUT5 #(
    .EQN("(~C*(D*~(E)*~((B*A))+D*E*~((B*A))+~(D)*E*(B*A)+D*E*(B*A)))"),
    .INIT(32'h0f080700))
    al_45894fd3 (
    .a(al_473186ca),
    .b(rx_clk_en),
    .c(al_ff9a7266),
    .d(al_c5bc3747),
    .e(al_a0f12bef[4]),
    .o(al_cb74bfe8));
  AL_DFF_X al_7239193 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_3252df70),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_9e8909aa));
  AL_DFF_X al_c62b6cf0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_6281ecee),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_8b7d9749));
  AL_DFF_0 al_3a13d081 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_7bec6b72),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9f0e53e2[0]));
  AL_DFF_0 al_7342e2e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_9f0e53e2[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9f0e53e2[1]));
  AL_DFF_0 al_9aa17f20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_9f0e53e2[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9f0e53e2[2]));
  AL_DFF_0 al_21f71d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_9f0e53e2[2]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9f0e53e2[3]));
  AL_DFF_0 al_85a86e23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_9f0e53e2[3]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9f0e53e2[4]));
  AL_DFF_0 al_d030be1b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_9f0e53e2[4]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9f0e53e2[5]));
  AL_DFF_0 al_8f915940 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f9cac200),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8867ef3c[0]));
  AL_DFF_0 al_5cd9f358 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_8867ef3c[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8867ef3c[1]));
  AL_DFF_0 al_70f44633 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_8867ef3c[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8867ef3c[2]));
  AL_DFF_0 al_76a0d527 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_d0a10128),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_628888c[0]));
  AL_DFF_0 al_a6cfd02c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_628888c[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_628888c[1]));
  AL_DFF_0 al_202cba8c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_628888c[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_628888c[2]));
  AL_DFF_0 al_8cab8790 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_628888c[2]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_628888c[3]));
  AL_DFF_X al_8c20c7a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_a0f12bef[1]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_316af0f0));
  AL_DFF_X al_cc463cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_6baf9e53),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_ce80051a));
  AL_DFF_X al_737f8928 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_2f3f17d),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_6ecd5054));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_8b97d87e (
    .a(rx_clk_en),
    .b(al_316af0f0),
    .o(al_15c18023));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    al_41f28a10 (
    .a(al_baa47a85),
    .b(al_b242ee60[0]),
    .c(al_db3c8a2c),
    .o(al_220ff640[0]));
  AL_MAP_LUT5 #(
    .EQN("(D@(C*(E@B@A)))"),
    .INIT(32'h6f909f60))
    al_87f26d42 (
    .a(al_27717189),
    .b(al_b242ee60[7]),
    .c(al_db3c8a2c),
    .d(al_39eeae1d[2]),
    .e(al_39eeae1d[24]),
    .o(al_220ff640[10]));
  AL_MAP_LUT6 #(
    .EQN("(E@(D*(F@C@B@A)))"),
    .INIT(64'h96ff690069ff9600))
    al_9037bcdb (
    .a(al_1c08f670),
    .b(al_fe465555),
    .c(al_b242ee60[7]),
    .d(al_db3c8a2c),
    .e(al_39eeae1d[3]),
    .f(al_39eeae1d[24]),
    .o(al_220ff640[11]));
  AL_MAP_LUT6 #(
    .EQN("(F@(E*(D@C@B@A)))"),
    .INIT(64'h9669ffff69960000))
    al_b33168c3 (
    .a(al_baa47a85),
    .b(al_bffbe171),
    .c(al_fe465555),
    .d(al_bb167cdd),
    .e(al_db3c8a2c),
    .f(al_39eeae1d[4]),
    .o(al_220ff640[12]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_b421560e (
    .a(al_b242ee60[5]),
    .b(al_39eeae1d[26]),
    .o(al_bb167cdd));
  AL_MAP_LUT4 #(
    .EQN("(D@C@B@A)"),
    .INIT(16'h6996))
    al_c1d27374 (
    .a(al_b242ee60[1]),
    .b(al_b242ee60[2]),
    .c(al_39eeae1d[29]),
    .d(al_39eeae1d[30]),
    .o(al_68c341e7));
  AL_MAP_LUT6 #(
    .EQN("(F@(E*(D@C@B@A)))"),
    .INIT(64'h9669ffff69960000))
    al_db345485 (
    .a(al_342f6170),
    .b(al_68c341e7),
    .c(al_3a7c57e3),
    .d(al_bb167cdd),
    .e(al_db3c8a2c),
    .f(al_39eeae1d[5]),
    .o(al_220ff640[13]));
  AL_MAP_LUT3 #(
    .EQN("(C@B@A)"),
    .INIT(8'h96))
    al_38af355c (
    .a(al_3a7c57e3),
    .b(al_b242ee60[3]),
    .c(al_39eeae1d[28]),
    .o(al_1c08f670));
  AL_MAP_LUT5 #(
    .EQN("(E@(D*~(C@B@A)))"),
    .INIT(32'h96ff6900))
    al_255637e7 (
    .a(al_5ea2be94[0]),
    .b(al_1c08f670),
    .c(al_bb167cdd),
    .d(al_db3c8a2c),
    .e(al_39eeae1d[6]),
    .o(al_220ff640[14]));
  AL_MAP_LUT5 #(
    .EQN("(E@(D*(C@B@A)))"),
    .INIT(32'h69ff9600))
    al_4636c9cd (
    .a(al_bffbe171),
    .b(al_3a7c57e3),
    .c(al_e3955cca),
    .d(al_db3c8a2c),
    .e(al_39eeae1d[7]),
    .o(al_220ff640[15]));
  AL_MAP_LUT5 #(
    .EQN("(D@(C*~(E@B@A)))"),
    .INIT(32'h9f606f90))
    al_18950224 (
    .a(al_bffbe171),
    .b(al_b242ee60[7]),
    .c(al_db3c8a2c),
    .d(al_39eeae1d[8]),
    .e(al_39eeae1d[24]),
    .o(al_220ff640[16]));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*~(B@A)))"),
    .INIT(16'h6f90))
    al_f0eb6bb4 (
    .a(al_68c341e7),
    .b(al_fe465555),
    .c(al_db3c8a2c),
    .d(al_39eeae1d[9]),
    .o(al_220ff640[17]));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*~(B@A)))"),
    .INIT(16'h6f90))
    al_f3c5b8e (
    .a(al_5ea2be94[0]),
    .b(al_bb167cdd),
    .c(al_db3c8a2c),
    .d(al_39eeae1d[10]),
    .o(al_220ff640[18]));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*(B@A)))"),
    .INIT(16'h9f60))
    al_ddb46ad0 (
    .a(al_3a7c57e3),
    .b(al_e3955cca),
    .c(al_db3c8a2c),
    .d(al_39eeae1d[11]),
    .o(al_220ff640[19]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    al_a05dbdb8 (
    .a(al_dacef8ff),
    .b(al_b242ee60[1]),
    .c(al_db3c8a2c),
    .o(al_220ff640[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(B*~(D@A)))"),
    .INIT(16'h78b4))
    al_eeb204fe (
    .a(al_b242ee60[3]),
    .b(al_db3c8a2c),
    .c(al_39eeae1d[12]),
    .d(al_39eeae1d[28]),
    .o(al_220ff640[20]));
  AL_MAP_LUT4 #(
    .EQN("(C@(B*~(D@A)))"),
    .INIT(16'h78b4))
    al_e70bbb7e (
    .a(al_b242ee60[2]),
    .b(al_db3c8a2c),
    .c(al_39eeae1d[13]),
    .d(al_39eeae1d[29]),
    .o(al_220ff640[21]));
  AL_MAP_LUT4 #(
    .EQN("(C@(B*~(D@A)))"),
    .INIT(16'h78b4))
    al_6e066b7b (
    .a(al_b242ee60[7]),
    .b(al_db3c8a2c),
    .c(al_39eeae1d[14]),
    .d(al_39eeae1d[24]),
    .o(al_220ff640[22]));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*~(B@A)))"),
    .INIT(16'h6f90))
    al_1ecc63dd (
    .a(al_baa47a85),
    .b(al_fe465555),
    .c(al_db3c8a2c),
    .d(al_39eeae1d[15]),
    .o(al_220ff640[23]));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*~(B@A)))"),
    .INIT(16'h6f90))
    al_4a693d91 (
    .a(al_342f6170),
    .b(al_bb167cdd),
    .c(al_db3c8a2c),
    .d(al_39eeae1d[16]),
    .o(al_220ff640[24]));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*(B@A)))"),
    .INIT(16'h9f60))
    al_e8db125a (
    .a(al_3a7c57e3),
    .b(al_bb167cdd),
    .c(al_db3c8a2c),
    .d(al_39eeae1d[17]),
    .o(al_220ff640[25]));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*(B@A)))"),
    .INIT(16'h9f60))
    al_a25f9240 (
    .a(al_1c08f670),
    .b(al_baa47a85),
    .c(al_db3c8a2c),
    .d(al_39eeae1d[18]),
    .o(al_220ff640[26]));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*(B@A)))"),
    .INIT(16'h9f60))
    al_272e586d (
    .a(al_342f6170),
    .b(al_bffbe171),
    .c(al_db3c8a2c),
    .d(al_39eeae1d[19]),
    .o(al_220ff640[27]));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*~(B@A)))"),
    .INIT(16'h6f90))
    al_161b3f16 (
    .a(al_68c341e7),
    .b(al_bb167cdd),
    .c(al_db3c8a2c),
    .d(al_39eeae1d[20]),
    .o(al_220ff640[28]));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*~(B@A)))"),
    .INIT(16'h6f90))
    al_dafd8e77 (
    .a(al_5ea2be94[0]),
    .b(al_3a7c57e3),
    .c(al_db3c8a2c),
    .d(al_39eeae1d[21]),
    .o(al_220ff640[29]));
  AL_MAP_LUT4 #(
    .EQN("(C*~((B@A))*~(D)+C*(B@A)*~(D)+~(C)*(B@A)*D+C*(B@A)*D)"),
    .INIT(16'h66f0))
    al_543c269a (
    .a(al_dacef8ff),
    .b(al_bb167cdd),
    .c(al_b242ee60[2]),
    .d(al_db3c8a2c),
    .o(al_220ff640[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(C*(E@B@A)))"),
    .INIT(32'h6f909f60))
    al_1e318be9 (
    .a(al_e3955cca),
    .b(al_b242ee60[3]),
    .c(al_db3c8a2c),
    .d(al_39eeae1d[22]),
    .e(al_39eeae1d[28]),
    .o(al_220ff640[30]));
  AL_MAP_LUT4 #(
    .EQN("(C@(B*~(D@A)))"),
    .INIT(16'h78b4))
    al_4a95e763 (
    .a(al_b242ee60[2]),
    .b(al_db3c8a2c),
    .c(al_39eeae1d[23]),
    .d(al_39eeae1d[29]),
    .o(al_220ff640[31]));
  AL_MAP_LUT5 #(
    .EQN("~(~D*~((C@B@A))*~(E)+~D*(C@B@A)*~(E)+~(~D)*(C@B@A)*E+~D*(C@B@A)*E)"),
    .INIT(32'h6969ff00))
    al_4ac73b68 (
    .a(al_342f6170),
    .b(al_3a7c57e3),
    .c(al_bb167cdd),
    .d(al_b242ee60[3]),
    .e(al_db3c8a2c),
    .o(al_220ff640[3]));
  AL_MAP_LUT5 #(
    .EQN("(D*~((C@B@A))*~(E)+D*(C@B@A)*~(E)+~(D)*(C@B@A)*E+D*(C@B@A)*E)"),
    .INIT(32'h9696ff00))
    al_1a5a18d4 (
    .a(al_1c08f670),
    .b(al_baa47a85),
    .c(al_bb167cdd),
    .d(al_b242ee60[4]),
    .e(al_db3c8a2c),
    .o(al_220ff640[4]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_e4a7ae41 (
    .a(al_b242ee60[4]),
    .b(al_39eeae1d[27]),
    .o(al_3a7c57e3));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_f2c313d (
    .a(al_342f6170),
    .b(al_baa47a85),
    .o(al_dacef8ff));
  AL_MAP_LUT5 #(
    .EQN("(D*~((C@B@A))*~(E)+D*(C@B@A)*~(E)+~(D)*(C@B@A)*E+D*(C@B@A)*E)"),
    .INIT(32'h9696ff00))
    al_3c059b6b (
    .a(al_dacef8ff),
    .b(al_bffbe171),
    .c(al_3a7c57e3),
    .d(al_b242ee60[5]),
    .e(al_db3c8a2c),
    .o(al_220ff640[5]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_611cce4e (
    .a(al_b242ee60[6]),
    .b(al_39eeae1d[25]),
    .o(al_fe465555));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_d7bd26ff (
    .a(al_b242ee60[0]),
    .b(al_39eeae1d[31]),
    .o(al_e3955cca));
  AL_MAP_LUT4 #(
    .EQN("(D@C@B@A)"),
    .INIT(16'h6996))
    al_bcf4c629 (
    .a(al_b242ee60[1]),
    .b(al_b242ee60[7]),
    .c(al_39eeae1d[24]),
    .d(al_39eeae1d[30]),
    .o(al_baa47a85));
  AL_MAP_LUT4 #(
    .EQN("(D@C@B@A)"),
    .INIT(16'h6996))
    al_e3d265a1 (
    .a(al_b242ee60[2]),
    .b(al_b242ee60[3]),
    .c(al_39eeae1d[28]),
    .d(al_39eeae1d[29]),
    .o(al_bffbe171));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_4ba3c754 (
    .a(al_fe465555),
    .b(al_e3955cca),
    .o(al_342f6170));
  AL_MAP_LUT3 #(
    .EQN("(C@B@A)"),
    .INIT(8'h96))
    al_2339bec9 (
    .a(al_e3955cca),
    .b(al_b242ee60[1]),
    .c(al_39eeae1d[30]),
    .o(al_5ea2be94[0]));
  AL_MAP_LUT6 #(
    .EQN("(D@(E*~(F@C@B@A)))"),
    .INIT(64'h6996ff009669ff00))
    al_dce79cdc (
    .a(al_5ea2be94[0]),
    .b(al_bffbe171),
    .c(al_bb167cdd),
    .d(al_b242ee60[6]),
    .e(al_db3c8a2c),
    .f(al_39eeae1d[25]),
    .o(al_220ff640[6]));
  AL_MAP_LUT4 #(
    .EQN("(D@C@B@A)"),
    .INIT(16'h6996))
    al_fc5940e (
    .a(al_3a7c57e3),
    .b(al_bb167cdd),
    .c(al_b242ee60[2]),
    .d(al_39eeae1d[29]),
    .o(al_27717189));
  AL_MAP_LUT5 #(
    .EQN("(C@(D*(E@B@A)))"),
    .INIT(32'h69f096f0))
    al_f5dad4a7 (
    .a(al_27717189),
    .b(al_e3955cca),
    .c(al_b242ee60[7]),
    .d(al_db3c8a2c),
    .e(al_39eeae1d[24]),
    .o(al_220ff640[7]));
  AL_MAP_LUT6 #(
    .EQN("(E@(D*(F@C@B@A)))"),
    .INIT(64'h96ff690069ff9600))
    al_a966b688 (
    .a(al_1c08f670),
    .b(al_fe465555),
    .c(al_b242ee60[7]),
    .d(al_db3c8a2c),
    .e(al_39eeae1d[0]),
    .f(al_39eeae1d[24]),
    .o(al_220ff640[8]));
  AL_MAP_LUT5 #(
    .EQN("(E@(D*(C@B@A)))"),
    .INIT(32'h69ff9600))
    al_d557ed68 (
    .a(al_bffbe171),
    .b(al_fe465555),
    .c(al_bb167cdd),
    .d(al_db3c8a2c),
    .e(al_39eeae1d[1]),
    .o(al_220ff640[9]));
  AL_DFF_X al_fd6d5ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_220ff640[0]),
    .en(al_15c18023),
    .sr(al_473186ca),
    .ss(1'b0),
    .q(al_39eeae1d[0]));
  AL_DFF_X al_c17312fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_220ff640[9]),
    .en(al_15c18023),
    .sr(al_473186ca),
    .ss(1'b0),
    .q(al_39eeae1d[9]));
  AL_DFF_X al_39618c84 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_220ff640[10]),
    .en(al_15c18023),
    .sr(al_473186ca),
    .ss(1'b0),
    .q(al_39eeae1d[10]));
  AL_DFF_X al_613c987f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_220ff640[11]),
    .en(al_15c18023),
    .sr(al_473186ca),
    .ss(1'b0),
    .q(al_39eeae1d[11]));
  AL_DFF_X al_227dd9f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_220ff640[12]),
    .en(al_15c18023),
    .sr(al_473186ca),
    .ss(1'b0),
    .q(al_39eeae1d[12]));
  AL_DFF_X al_66db8d6c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_220ff640[13]),
    .en(al_15c18023),
    .sr(al_473186ca),
    .ss(1'b0),
    .q(al_39eeae1d[13]));
  AL_DFF_X al_affeee8c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_220ff640[14]),
    .en(al_15c18023),
    .sr(al_473186ca),
    .ss(1'b0),
    .q(al_39eeae1d[14]));
  AL_DFF_X al_8f6374a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_220ff640[15]),
    .en(al_15c18023),
    .sr(al_473186ca),
    .ss(1'b0),
    .q(al_39eeae1d[15]));
  AL_DFF_X al_31789fa7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_220ff640[16]),
    .en(al_15c18023),
    .sr(al_473186ca),
    .ss(1'b0),
    .q(al_39eeae1d[16]));
  AL_DFF_X al_4c6c544b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_220ff640[17]),
    .en(al_15c18023),
    .sr(al_473186ca),
    .ss(1'b0),
    .q(al_39eeae1d[17]));
  AL_DFF_X al_f8a67a68 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_220ff640[18]),
    .en(al_15c18023),
    .sr(al_473186ca),
    .ss(1'b0),
    .q(al_39eeae1d[18]));
  AL_DFF_X al_4e48ffef (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_220ff640[1]),
    .en(al_15c18023),
    .sr(al_473186ca),
    .ss(1'b0),
    .q(al_39eeae1d[1]));
  AL_DFF_X al_a4df6c7f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_220ff640[19]),
    .en(al_15c18023),
    .sr(al_473186ca),
    .ss(1'b0),
    .q(al_39eeae1d[19]));
  AL_DFF_X al_70146b96 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_220ff640[20]),
    .en(al_15c18023),
    .sr(al_473186ca),
    .ss(1'b0),
    .q(al_39eeae1d[20]));
  AL_DFF_X al_2bf60cfe (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_220ff640[21]),
    .en(al_15c18023),
    .sr(al_473186ca),
    .ss(1'b0),
    .q(al_39eeae1d[21]));
  AL_DFF_X al_8f704f41 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_220ff640[22]),
    .en(al_15c18023),
    .sr(al_473186ca),
    .ss(1'b0),
    .q(al_39eeae1d[22]));
  AL_DFF_X al_33c809d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_220ff640[23]),
    .en(al_15c18023),
    .sr(al_473186ca),
    .ss(1'b0),
    .q(al_39eeae1d[23]));
  AL_DFF_X al_dbc8358a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_220ff640[24]),
    .en(al_15c18023),
    .sr(al_473186ca),
    .ss(1'b0),
    .q(al_39eeae1d[24]));
  AL_DFF_X al_c33646d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_220ff640[25]),
    .en(al_15c18023),
    .sr(al_473186ca),
    .ss(1'b0),
    .q(al_39eeae1d[25]));
  AL_DFF_X al_9542fc4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_220ff640[26]),
    .en(al_15c18023),
    .sr(al_473186ca),
    .ss(1'b0),
    .q(al_39eeae1d[26]));
  AL_DFF_X al_8645f0e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_220ff640[27]),
    .en(al_15c18023),
    .sr(al_473186ca),
    .ss(1'b0),
    .q(al_39eeae1d[27]));
  AL_DFF_X al_1bf9628c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_220ff640[28]),
    .en(al_15c18023),
    .sr(al_473186ca),
    .ss(1'b0),
    .q(al_39eeae1d[28]));
  AL_DFF_X al_8cb0b987 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_220ff640[2]),
    .en(al_15c18023),
    .sr(al_473186ca),
    .ss(1'b0),
    .q(al_39eeae1d[2]));
  AL_DFF_X al_b0a3a642 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_220ff640[29]),
    .en(al_15c18023),
    .sr(al_473186ca),
    .ss(1'b0),
    .q(al_39eeae1d[29]));
  AL_DFF_X al_332aad13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_220ff640[30]),
    .en(al_15c18023),
    .sr(al_473186ca),
    .ss(1'b0),
    .q(al_39eeae1d[30]));
  AL_DFF_X al_f3b1fd7e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_220ff640[31]),
    .en(al_15c18023),
    .sr(al_473186ca),
    .ss(1'b0),
    .q(al_39eeae1d[31]));
  AL_DFF_X al_1b6fba9d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_220ff640[3]),
    .en(al_15c18023),
    .sr(al_473186ca),
    .ss(1'b0),
    .q(al_39eeae1d[3]));
  AL_DFF_X al_9fbf18f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_220ff640[4]),
    .en(al_15c18023),
    .sr(al_473186ca),
    .ss(1'b0),
    .q(al_39eeae1d[4]));
  AL_DFF_X al_725f362 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_220ff640[5]),
    .en(al_15c18023),
    .sr(al_473186ca),
    .ss(1'b0),
    .q(al_39eeae1d[5]));
  AL_DFF_X al_d59d370c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_220ff640[6]),
    .en(al_15c18023),
    .sr(al_473186ca),
    .ss(1'b0),
    .q(al_39eeae1d[6]));
  AL_DFF_X al_967b3f63 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_220ff640[7]),
    .en(al_15c18023),
    .sr(al_473186ca),
    .ss(1'b0),
    .q(al_39eeae1d[7]));
  AL_DFF_X al_728bd1f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_220ff640[8]),
    .en(al_15c18023),
    .sr(al_473186ca),
    .ss(1'b0),
    .q(al_39eeae1d[8]));
  AL_DFF_X al_7a5976fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_c5c11e98),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_af3abf3a));
  AL_DFF_X al_e49140c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1217cf69),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_a14eea73));
  AL_DFF_X al_862a74b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_164531d8),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_fa54303d));
  AL_DFF_X al_cc73b023 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_88b7c5fc),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_e4bdca8a));
  AL_DFF_X al_323dcfc0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1bae0f4e),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_c8fffdaf));
  AL_DFF_X al_8f181c69 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_535d21bf),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_1c648f36));
  AL_DFF_X al_2fea96b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_6a75b886),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_8aec7267));
  AL_DFF_X al_7b6bbdee (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_4529840c),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_1af0ad5e));
  AL_DFF_X al_e717b2b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_7f95b06f),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_a1ace55b));
  AL_DFF_X al_6c531e03 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_db02221b),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_cd9c4b15));
  AL_DFF_X al_22eed131 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_bbb4d320),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_8769457b));
  AL_DFF_X al_26980342 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_33991d35),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(al_ff9a7266),
    .q(al_31732ee5));
  AL_DFF_X al_f39590c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_fdcd79c7),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_32839ce1));
  AL_DFF_X al_aee1d3b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_3714f7a3),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_e3b877ad));
  AL_DFF_X al_5af58cdc (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_506bb8a),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_75c3c1c0));
  AL_DFF_X al_560ce7e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e3b877ad),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_dc6fb7d9));
  AL_DFF_X al_955457b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_6333de40),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_e1d5aa87));
  AL_DFF_X al_c65592c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_aa43251),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_6c890ee8));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*~(C*B)))"),
    .INIT(16'h5540))
    al_6b8295f8 (
    .a(al_9907ae47),
    .b(al_77df94be),
    .c(al_75c3c1c0),
    .d(al_c8fffdaf),
    .o(al_1bae0f4e));
  AL_MAP_LUT5 #(
    .EQN("(~C*~B*~A*~(E@D))"),
    .INIT(32'h01000001))
    al_cf1851e4 (
    .a(al_3a7c57e3),
    .b(al_fe465555),
    .c(al_bb167cdd),
    .d(al_b242ee60[1]),
    .e(al_39eeae1d[30]),
    .o(al_20c70ab1));
  AL_MAP_LUT6 #(
    .EQN("(~B*A*~(E@D)*~(F@C))"),
    .INIT(64'h2000002002000002))
    al_454a2094 (
    .a(al_20c70ab1),
    .b(al_e3955cca),
    .c(al_b242ee60[2]),
    .d(al_b242ee60[7]),
    .e(al_39eeae1d[24]),
    .f(al_39eeae1d[29]),
    .o(al_458cb894));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D@B)))"),
    .INIT(16'h70d0))
    al_d1307868 (
    .a(al_458cb894),
    .b(al_b242ee60[3]),
    .c(al_e06bfe23),
    .d(al_39eeae1d[28]),
    .o(al_164531d8));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_6619a508 (
    .a(al_c2569e9f),
    .b(al_db0897ce),
    .c(al_7701781b),
    .o(al_8cf1eeca));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(~B*~A*~(E*~C)))"),
    .INIT(32'h00ef00ee))
    al_e54ea671 (
    .a(al_8cf1eeca),
    .b(al_88b7c5fc),
    .c(al_ce80051a),
    .d(al_9907ae47),
    .e(al_535d21bf),
    .o(al_6a75b886));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~D*~C*~A))"),
    .INIT(16'h3332))
    al_820054e7 (
    .a(al_e2923d0b),
    .b(al_9907ae47),
    .c(al_af3abf3a),
    .d(al_4df60ad5),
    .o(al_c5c11e98));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_448fe178 (
    .a(al_fa54303d),
    .b(al_8aec7267),
    .o(al_88b7c5fc));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_9fe573d5 (
    .a(al_9907ae47),
    .b(al_31732ee5),
    .o(al_aa43251));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*~A)"),
    .INIT(32'h00000004))
    al_eeffab7a (
    .a(al_88b7c5fc),
    .b(al_aa43251),
    .c(al_a1ace55b),
    .d(al_e3b877ad),
    .e(al_e1d5aa87),
    .o(al_db02221b));
  AL_MAP_LUT5 #(
    .EQN("(B*~(~E*~D*~C*~A))"),
    .INIT(32'hccccccc8))
    al_96baf562 (
    .a(al_88b7c5fc),
    .b(al_aa43251),
    .c(al_a1ace55b),
    .d(al_e3b877ad),
    .e(al_e1d5aa87),
    .o(al_1217cf69));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_282469c1 (
    .a(al_cca5b6a5),
    .b(al_a1ace55b),
    .o(al_fdcd79c7));
  AL_MAP_LUT6 #(
    .EQN("(~(~F*E)*~(~(D*~B)*~(C*~A)))"),
    .INIT(64'h7350735000007350))
    al_407943f6 (
    .a(al_d632949b),
    .b(al_cc4e6731),
    .c(al_d0ecc99e),
    .d(al_8e811a01),
    .e(al_75c3c1c0),
    .f(al_c8fffdaf),
    .o(al_83c2aae7));
  AL_MAP_LUT6 #(
    .EQN("(C*~(~A*~(~F*~E*~D*~B)))"),
    .INIT(64'ha0a0a0a0a0a0a0b0))
    al_cfc4e36a (
    .a(al_83c2aae7),
    .b(al_d632949b),
    .c(al_2ff03e70),
    .d(al_994b00c4),
    .e(al_d0ecc99e),
    .f(al_cca5b6a5),
    .o(al_1adec7e7));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(~E*~A*~(~D*C)))"),
    .INIT(32'h33332232))
    al_2ebf403d (
    .a(al_1adec7e7),
    .b(al_9907ae47),
    .c(al_e06bfe23),
    .d(al_c8fffdaf),
    .e(al_a1ace55b),
    .o(al_7f95b06f));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    al_61da6c32 (
    .a(al_473186ca),
    .b(al_9907ae47),
    .c(al_31732ee5),
    .o(al_33991d35));
  AL_MAP_LUT6 #(
    .EQN("(E*~D*~C*~A*~(F*~B))"),
    .INIT(64'h0004000000050000))
    al_8d273963 (
    .a(al_535d21bf),
    .b(al_aac09418[2]),
    .c(al_aac09418[3]),
    .d(al_aac09418[9]),
    .e(al_aac09418[10]),
    .f(al_391ec013),
    .o(al_23cb1fcc));
  AL_MAP_LUT6 #(
    .EQN("(~F*~(~E*D*~C*B*A))"),
    .INIT(64'h00000000fffff7ff))
    al_8b1dc2d7 (
    .a(al_23cb1fcc),
    .b(al_7557c0dc),
    .c(al_aac09418[0]),
    .d(al_aac09418[1]),
    .e(al_aac09418[4]),
    .f(al_e3b877ad),
    .o(al_407365eb));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_2cff9c73 (
    .a(al_407365eb),
    .b(al_ff67665e),
    .c(al_9907ae47),
    .o(al_3714f7a3));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*B*A)"),
    .INIT(32'h00000080))
    al_ace9ad92 (
    .a(al_aac09418[2]),
    .b(al_aac09418[3]),
    .c(al_aac09418[5]),
    .d(al_aac09418[6]),
    .e(al_aac09418[7]),
    .o(al_1973de82));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    al_71978725 (
    .a(al_1973de82),
    .b(al_aac09418[0]),
    .c(al_aac09418[1]),
    .d(al_aac09418[4]),
    .o(al_506bb8a));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C@B))"),
    .INIT(8'hbe))
    al_861bf94a (
    .a(al_76ee0125),
    .b(al_bcf9a5e2),
    .c(al_be957c85[0]),
    .o(al_1ac19429[0]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D@(C*B)))"),
    .INIT(16'h1540))
    al_a51ecd2a (
    .a(al_76ee0125),
    .b(al_bcf9a5e2),
    .c(al_be957c85[0]),
    .d(al_be957c85[1]),
    .o(al_1ac19429[1]));
  AL_MAP_LUT5 #(
    .EQN("(~A*(E@(D*C*B)))"),
    .INIT(32'h15554000))
    al_d5b5ca20 (
    .a(al_76ee0125),
    .b(al_bcf9a5e2),
    .c(al_be957c85[0]),
    .d(al_be957c85[1]),
    .e(al_be957c85[2]),
    .o(al_1ac19429[2]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D@(C*B)))"),
    .INIT(16'h1540))
    al_c8fe9b35 (
    .a(al_76ee0125),
    .b(al_bcf9a5e2),
    .c(al_8999d24b),
    .d(al_be957c85[3]),
    .o(al_1ac19429[3]));
  AL_MAP_LUT3 #(
    .EQN("(~A*(C@B))"),
    .INIT(8'h14))
    al_1e5c5601 (
    .a(al_76ee0125),
    .b(al_1629ae4d),
    .c(al_be957c85[4]),
    .o(al_1ac19429[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_7b8f54e4 (
    .a(al_bcf9a5e2),
    .b(al_8999d24b),
    .c(al_be957c85[3]),
    .o(al_1629ae4d));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D@(C*B)))"),
    .INIT(16'h1540))
    al_93a71a89 (
    .a(al_76ee0125),
    .b(al_1629ae4d),
    .c(al_be957c85[4]),
    .d(al_be957c85[5]),
    .o(al_1ac19429[5]));
  AL_MAP_LUT3 #(
    .EQN("(~A*(C@B))"),
    .INIT(8'h14))
    al_6edb05f7 (
    .a(al_76ee0125),
    .b(al_3e13fa86),
    .c(al_be957c85[6]),
    .o(al_1ac19429[6]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D@(C*B)))"),
    .INIT(16'h1540))
    al_88032ada (
    .a(al_76ee0125),
    .b(al_3e13fa86),
    .c(al_be957c85[6]),
    .d(al_be957c85[7]),
    .o(al_1ac19429[7]));
  AL_MAP_LUT5 #(
    .EQN("(~A*(E@(D*C*B)))"),
    .INIT(32'h15554000))
    al_eeabed09 (
    .a(al_76ee0125),
    .b(al_3e13fa86),
    .c(al_be957c85[6]),
    .d(al_be957c85[7]),
    .e(al_be957c85[8]),
    .o(al_1ac19429[8]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    al_d00ac00 (
    .a(al_6cdf2816),
    .b(al_7701781b),
    .c(al_d5b2f5c4),
    .d(al_614db0a6),
    .o(al_bbb4d320));
  AL_MAP_LUT6 #(
    .EQN("(~A*~(~F*~(E*D*C*B)))"),
    .INIT(64'h5555555540000000))
    al_4d4b7e16 (
    .a(al_76ee0125),
    .b(al_3e13fa86),
    .c(al_be957c85[6]),
    .d(al_be957c85[7]),
    .e(al_be957c85[8]),
    .f(al_be957c85[9]),
    .o(al_1ac19429[9]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_5c07630f (
    .a(al_bbb4d320),
    .b(al_8769457b),
    .o(al_76ee0125));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_6fee958 (
    .a(al_49bc5cf4),
    .b(al_be957c85[6]),
    .c(al_be957c85[9]),
    .o(al_aeadc72a));
  AL_MAP_LUT6 #(
    .EQN("(~B*~(~E*~D*A*~(~F*C)))"),
    .INIT(64'h3333331133333331))
    al_834fd92c (
    .a(al_6cdf2816),
    .b(al_aeadc72a),
    .c(al_7701781b),
    .d(al_d5b2f5c4),
    .e(al_614db0a6),
    .f(al_1af0ad5e),
    .o(al_bcf9a5e2));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_b80d1671 (
    .a(al_be957c85[0]),
    .b(al_be957c85[1]),
    .c(al_be957c85[2]),
    .o(al_8999d24b));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    al_2612bf54 (
    .a(al_bcf9a5e2),
    .b(al_8999d24b),
    .c(al_be957c85[3]),
    .d(al_be957c85[4]),
    .e(al_be957c85[5]),
    .o(al_3e13fa86));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(D*~(C*B)))"),
    .INIT(16'hbfaa))
    al_b577922e (
    .a(al_76ee0125),
    .b(al_7701781b),
    .c(al_1c648f36),
    .d(al_1af0ad5e),
    .o(al_4529840c));
  AL_MAP_LUT6 #(
    .EQN("(F*~(E*B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A)))"),
    .INIT(64'h3b7fffff00000000))
    al_8e45305f (
    .a(al_49bc5cf4),
    .b(al_7701781b),
    .c(al_aea26701[6]),
    .d(al_aea26701[9]),
    .e(al_1c648f36),
    .f(al_e1d5aa87),
    .o(al_d8bfe065));
  AL_MAP_LUT6 #(
    .EQN("((B*~(F*~E*C))*~(D)*~(A)+(B*~(F*~E*C))*D*~(A)+~((B*~(F*~E*C)))*D*A+(B*~(F*~E*C))*D*A)"),
    .INIT(64'hee44ae04ee44ee44))
    al_d14f00ff (
    .a(al_76ee0125),
    .b(al_d8bfe065),
    .c(al_aeadc72a),
    .d(al_54d691ed),
    .e(al_7701781b),
    .f(al_1af0ad5e),
    .o(al_6333de40));
  AL_DFF_X al_9ffc6f9f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1ac19429[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(al_ff9a7266),
    .q(al_be957c85[0]));
  AL_DFF_X al_4d9128ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1ac19429[9]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_be957c85[9]));
  AL_DFF_X al_fafbf17d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1ac19429[1]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_be957c85[1]));
  AL_DFF_X al_be2afad5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1ac19429[2]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_be957c85[2]));
  AL_DFF_X al_852c4583 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1ac19429[3]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_be957c85[3]));
  AL_DFF_X al_787b34c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1ac19429[4]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_be957c85[4]));
  AL_DFF_X al_86f1ba10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1ac19429[5]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_be957c85[5]));
  AL_DFF_X al_d43f759a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1ac19429[6]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_be957c85[6]));
  AL_DFF_X al_4059679b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1ac19429[7]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_be957c85[7]));
  AL_DFF_X al_317123aa (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1ac19429[8]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_be957c85[8]));
  AL_DFF_X al_2433e00b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_be957c85[9]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_aea26701[9]));
  AL_DFF_X al_6813e772 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_be957c85[6]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_aea26701[6]));
  AL_DFF_X al_ddc3d729 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_27161c58),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_823fecd4));
  AL_DFF_X al_c16a0462 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_823fecd4),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_1180f8c0));
  AL_DFF_X al_5dd703ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1180f8c0),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_8b780845));
  AL_DFF_X al_e38a1f28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f7483e6d),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_735aa681));
  AL_DFF_X al_a2c4ff88 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_735aa681),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_8e811a01));
  AL_DFF_X al_e51337de (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_949a133d),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_4f1a9685));
  AL_DFF_X al_590dc1e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_a0088870),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_db3c8a2c));
  AL_DFF_X al_9293083a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_4cf5bca0),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_2c7a1247));
  AL_DFF_X al_1626a421 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_a396e89f),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_cac2565f));
  AL_DFF_X al_5d690016 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e1409b5e),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_fe00f314));
  AL_DFF_X al_34582806 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_18337cf7),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_994b00c4));
  AL_DFF_X al_36a0d24a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0947bb5),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_1ed21a96));
  AL_DFF_X al_d65767b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_8996909b),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_51ab8bb8));
  AL_DFF_X al_8008ec9d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_618737cb),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_a783ebfd));
  AL_DFF_X al_f1e30d9a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_4f9f38e2),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_ed990b15));
  AL_DFF_X al_ba3c2fef (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_34aaf187),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_4f9f38e2));
  AL_DFF_X al_59f2d056 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_38b760cc),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d0ecc99e));
  AL_MAP_LUT6 #(
    .EQN("(~C*(A*B*~((E*D))*~(F)+A*B*(E*D)*~(F)+~(A)*~(B)*~((E*D))*F+A*~(B)*~((E*D))*F+~(A)*B*~((E*D))*F+A*B*~((E*D))*F+~(A)*~(B)*(E*D)*F+A*~(B)*(E*D)*F+A*B*(E*D)*F))"),
    .INIT(64'h0b0f0f0f08080808))
    al_e0be8722 (
    .a(al_31ba2088),
    .b(rx_clk_en),
    .c(al_ff9a7266),
    .d(al_2e8ff7ab),
    .e(al_54f03dbf[1]),
    .f(al_d0ecc99e),
    .o(al_38b760cc));
  AL_MAP_LUT5 #(
    .EQN("(E*~(~D*~(C*B*A)))"),
    .INIT(32'hff800000))
    al_878ff298 (
    .a(al_b242ee60[1]),
    .b(al_b242ee60[2]),
    .c(al_b242ee60[3]),
    .d(al_b242ee60[4]),
    .e(al_b242ee60[5]),
    .o(al_7c0134d3));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*~C*~B*~A)"),
    .INIT(64'h0100000000000000))
    al_e6ba0525 (
    .a(al_7c0134d3),
    .b(al_b242ee60[6]),
    .c(al_b242ee60[7]),
    .d(al_2e8ff7ab),
    .e(al_54f03dbf[1]),
    .f(al_a783ebfd),
    .o(al_31ba2088));
  AL_DFF_X al_8bc5a625 (
    .ar(al_ff9a7266),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_c2569e9f),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccf401cd));
  AL_DFF_X al_c271bc99 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_63101725),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(al_ff9a7266),
    .q(al_cca5b6a5));
  AL_DFF_X al_40718249 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_d6a2be89[1]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_391ec013));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_7b5c85af (
    .a(1'b0),
    .o({al_25b9a235,open_n6}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_1d1635f3 (
    .a(al_cbc62139[0]),
    .b(1'b1),
    .c(al_25b9a235),
    .o({al_c9d3334,al_c86ca47d[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ef6071dc (
    .a(al_cbc62139[1]),
    .b(1'b0),
    .c(al_c9d3334),
    .o({al_a021098c,al_c86ca47d[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_6cccdfc5 (
    .a(al_cbc62139[2]),
    .b(1'b0),
    .c(al_a021098c),
    .o({al_e0f968c1,al_c86ca47d[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f8ba1dad (
    .a(al_cbc62139[3]),
    .b(1'b0),
    .c(al_e0f968c1),
    .o({al_40bf3e87,al_c86ca47d[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_11445499 (
    .a(al_cbc62139[4]),
    .b(1'b0),
    .c(al_40bf3e87),
    .o({al_baff81fb,al_c86ca47d[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_5c040c8c (
    .a(al_cbc62139[5]),
    .b(1'b0),
    .c(al_baff81fb),
    .o({al_e44d618,al_c86ca47d[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a673b89b (
    .a(al_cbc62139[6]),
    .b(1'b0),
    .c(al_e44d618),
    .o({al_6ab58fb5,al_c86ca47d[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_9c2773a4 (
    .a(al_cbc62139[7]),
    .b(1'b0),
    .c(al_6ab58fb5),
    .o({al_37c809df,al_c86ca47d[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e32ad97a (
    .a(al_cbc62139[8]),
    .b(1'b0),
    .c(al_37c809df),
    .o({al_1d552e04,al_c86ca47d[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_69c1249e (
    .a(al_cbc62139[9]),
    .b(1'b0),
    .c(al_1d552e04),
    .o({al_307af410,al_c86ca47d[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_552d4d8c (
    .a(al_cbc62139[10]),
    .b(1'b0),
    .c(al_307af410),
    .o({al_1e561c50,al_c86ca47d[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_8e8a9fb (
    .a(al_cbc62139[11]),
    .b(1'b0),
    .c(al_1e561c50),
    .o({al_9b855829,al_c86ca47d[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_7e9f6953 (
    .a(al_cbc62139[12]),
    .b(1'b0),
    .c(al_9b855829),
    .o({al_41381f51,al_c86ca47d[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ec838b5f (
    .a(al_cbc62139[13]),
    .b(1'b0),
    .c(al_41381f51),
    .o({al_2e700a59,al_c86ca47d[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a9d54d64 (
    .a(al_cbc62139[14]),
    .b(1'b0),
    .c(al_2e700a59),
    .o({open_n7,al_c86ca47d[14]}));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    al_7c0aa89d (
    .a(rx_clk_en),
    .b(al_cbc62139[14]),
    .c(al_ccf401cd),
    .o(al_e7a9a14d));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .INIT(16'h4540))
    al_f9f8fff (
    .a(al_473186ca),
    .b(al_cbc62139[0]),
    .c(al_cbc62139[14]),
    .d(al_c86ca47d[0]),
    .o(al_92477e6d[0]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .INIT(16'h4540))
    al_aa281eac (
    .a(al_473186ca),
    .b(al_cbc62139[10]),
    .c(al_cbc62139[14]),
    .d(al_c86ca47d[10]),
    .o(al_92477e6d[10]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .INIT(16'h4540))
    al_c66eb31c (
    .a(al_473186ca),
    .b(al_cbc62139[11]),
    .c(al_cbc62139[14]),
    .d(al_c86ca47d[11]),
    .o(al_92477e6d[11]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .INIT(16'h4540))
    al_fe5c4da9 (
    .a(al_473186ca),
    .b(al_cbc62139[12]),
    .c(al_cbc62139[14]),
    .d(al_c86ca47d[12]),
    .o(al_92477e6d[12]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .INIT(16'h4540))
    al_930ecf3b (
    .a(al_473186ca),
    .b(al_cbc62139[13]),
    .c(al_cbc62139[14]),
    .d(al_c86ca47d[13]),
    .o(al_92477e6d[13]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    al_a33ca611 (
    .a(al_473186ca),
    .b(al_cbc62139[14]),
    .c(al_c86ca47d[14]),
    .o(al_92477e6d[14]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .INIT(16'h4540))
    al_d834f745 (
    .a(al_473186ca),
    .b(al_cbc62139[1]),
    .c(al_cbc62139[14]),
    .d(al_c86ca47d[1]),
    .o(al_92477e6d[1]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .INIT(16'h4540))
    al_76e839c9 (
    .a(al_473186ca),
    .b(al_cbc62139[2]),
    .c(al_cbc62139[14]),
    .d(al_c86ca47d[2]),
    .o(al_92477e6d[2]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .INIT(16'h4540))
    al_14ed2af1 (
    .a(al_473186ca),
    .b(al_cbc62139[3]),
    .c(al_cbc62139[14]),
    .d(al_c86ca47d[3]),
    .o(al_92477e6d[3]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .INIT(16'h4540))
    al_b90108ff (
    .a(al_473186ca),
    .b(al_cbc62139[4]),
    .c(al_cbc62139[14]),
    .d(al_c86ca47d[4]),
    .o(al_92477e6d[4]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .INIT(16'h4540))
    al_e4d98d34 (
    .a(al_473186ca),
    .b(al_cbc62139[5]),
    .c(al_cbc62139[14]),
    .d(al_c86ca47d[5]),
    .o(al_92477e6d[5]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .INIT(16'h4540))
    al_9afa2f5a (
    .a(al_473186ca),
    .b(al_cbc62139[6]),
    .c(al_cbc62139[14]),
    .d(al_c86ca47d[6]),
    .o(al_92477e6d[6]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .INIT(16'h4540))
    al_a0560213 (
    .a(al_473186ca),
    .b(al_cbc62139[7]),
    .c(al_cbc62139[14]),
    .d(al_c86ca47d[7]),
    .o(al_92477e6d[7]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .INIT(16'h4540))
    al_e38e4950 (
    .a(al_473186ca),
    .b(al_cbc62139[8]),
    .c(al_cbc62139[14]),
    .d(al_c86ca47d[8]),
    .o(al_92477e6d[8]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .INIT(16'h4540))
    al_ea4b0aa0 (
    .a(al_473186ca),
    .b(al_cbc62139[9]),
    .c(al_cbc62139[14]),
    .d(al_c86ca47d[9]),
    .o(al_92477e6d[9]));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    al_5a8105e (
    .a(al_d5b2f5c4),
    .b(al_e06bfe23),
    .c(al_54f03dbf[0]),
    .d(al_2ff03e70),
    .o(al_e4f71d03));
  AL_MAP_LUT5 #(
    .EQN("((~E*D*~C)*~(B)*~(A)+(~E*D*~C)*B*~(A)+~((~E*D*~C))*B*A+(~E*D*~C)*B*A)"),
    .INIT(32'h88888d88))
    al_638d2447 (
    .a(al_e4f71d03),
    .b(al_b242ee60[0]),
    .c(al_9907ae47),
    .d(al_4f9f38e2),
    .e(al_7bec6b72),
    .o(al_34aaf187));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(E*~(B)*~((D*C))+E*B*~((D*C))+~(E)*B*(D*C)+E*B*(D*C)))"),
    .INIT(32'hefffeaaa))
    al_5620a6c7 (
    .a(al_473186ca),
    .b(al_b242ee60[0]),
    .c(al_2e8ff7ab),
    .d(al_54f03dbf[1]),
    .e(al_14016c23[0]),
    .o(al_f0afd253[0]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'hfbea))
    al_c4734e63 (
    .a(al_473186ca),
    .b(al_d1451a79),
    .c(al_b242ee60[2]),
    .d(al_14016c23[10]),
    .o(al_f0afd253[10]));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(E*~(B)*~((D*C))+E*B*~((D*C))+~(E)*B*(D*C)+E*B*(D*C)))"),
    .INIT(32'hefffeaaa))
    al_40f9af81 (
    .a(al_473186ca),
    .b(al_b242ee60[1]),
    .c(al_2e8ff7ab),
    .d(al_54f03dbf[1]),
    .e(al_14016c23[1]),
    .o(al_f0afd253[1]));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(E*~(B)*~((D*C))+E*B*~((D*C))+~(E)*B*(D*C)+E*B*(D*C)))"),
    .INIT(32'hefffeaaa))
    al_5f04589a (
    .a(al_473186ca),
    .b(al_b242ee60[2]),
    .c(al_2e8ff7ab),
    .d(al_54f03dbf[1]),
    .e(al_14016c23[2]),
    .o(al_f0afd253[2]));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(E*~(B)*~((D*C))+E*B*~((D*C))+~(E)*B*(D*C)+E*B*(D*C)))"),
    .INIT(32'hefffeaaa))
    al_5bd722e8 (
    .a(al_473186ca),
    .b(al_b242ee60[3]),
    .c(al_2e8ff7ab),
    .d(al_54f03dbf[1]),
    .e(al_14016c23[3]),
    .o(al_f0afd253[3]));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(E*~(B)*~((D*C))+E*B*~((D*C))+~(E)*B*(D*C)+E*B*(D*C)))"),
    .INIT(32'hefffeaaa))
    al_6b026c37 (
    .a(al_473186ca),
    .b(al_b242ee60[4]),
    .c(al_2e8ff7ab),
    .d(al_54f03dbf[1]),
    .e(al_14016c23[4]),
    .o(al_f0afd253[4]));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(E*~(B)*~((D*C))+E*B*~((D*C))+~(E)*B*(D*C)+E*B*(D*C)))"),
    .INIT(32'hefffeaaa))
    al_30ee9861 (
    .a(al_473186ca),
    .b(al_b242ee60[5]),
    .c(al_2e8ff7ab),
    .d(al_54f03dbf[1]),
    .e(al_14016c23[5]),
    .o(al_f0afd253[5]));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(E*~(B)*~((D*C))+E*B*~((D*C))+~(E)*B*(D*C)+E*B*(D*C)))"),
    .INIT(32'hefffeaaa))
    al_f94741b4 (
    .a(al_473186ca),
    .b(al_b242ee60[6]),
    .c(al_2e8ff7ab),
    .d(al_54f03dbf[1]),
    .e(al_14016c23[6]),
    .o(al_f0afd253[6]));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(E*~(B)*~((D*C))+E*B*~((D*C))+~(E)*B*(D*C)+E*B*(D*C)))"),
    .INIT(32'hefffeaaa))
    al_1e5b79f3 (
    .a(al_473186ca),
    .b(al_b242ee60[7]),
    .c(al_2e8ff7ab),
    .d(al_54f03dbf[1]),
    .e(al_14016c23[7]),
    .o(al_f0afd253[7]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'hfbea))
    al_a66e98eb (
    .a(al_473186ca),
    .b(al_d1451a79),
    .c(al_b242ee60[0]),
    .d(al_14016c23[8]),
    .o(al_f0afd253[8]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'hfbea))
    al_9f8990ee (
    .a(al_473186ca),
    .b(al_d1451a79),
    .c(al_b242ee60[1]),
    .d(al_14016c23[9]),
    .o(al_f0afd253[9]));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*~B*A)"),
    .INIT(32'h00020000))
    al_6d7059a0 (
    .a(al_d1451a79),
    .b(al_b242ee60[4]),
    .c(al_b242ee60[5]),
    .d(al_b242ee60[6]),
    .e(al_b242ee60[7]),
    .o(al_6ec43dd2));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*C*B*A)"),
    .INIT(64'h0000000000000080))
    al_fc603e98 (
    .a(al_6ec43dd2),
    .b(al_531e5772),
    .c(al_b242ee60[0]),
    .d(al_b242ee60[1]),
    .e(al_b242ee60[2]),
    .f(al_b242ee60[3]),
    .o(al_87b441ee));
  AL_MAP_LUT6 #(
    .EQN("((F*~B)*~((E*A))*~((D*C))+(F*~B)*(E*A)*~((D*C))+~((F*~B))*(E*A)*(D*C)+(F*~B)*(E*A)*(D*C))"),
    .INIT(64'ha3330333a0000000))
    al_9b2d0539 (
    .a(al_d86c9f70),
    .b(al_9907ae47),
    .c(al_2e8ff7ab),
    .d(al_54f03dbf[1]),
    .e(al_d6a2be89[0]),
    .f(al_d6a2be89[1]),
    .o(al_59c37d06));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    al_a33ed433 (
    .a(al_b242ee60[0]),
    .b(al_b242ee60[1]),
    .c(al_b242ee60[2]),
    .d(al_b242ee60[3]),
    .o(al_1ff7640d));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    al_12eed2b2 (
    .a(al_1ff7640d),
    .b(al_b242ee60[4]),
    .c(al_b242ee60[5]),
    .d(al_b242ee60[6]),
    .e(al_b242ee60[7]),
    .o(al_cc14f446));
  AL_MAP_LUT6 #(
    .EQN("((F*~B)*~((E*A))*~((D*C))+(F*~B)*(E*A)*~((D*C))+~((F*~B))*(E*A)*(D*C)+(F*~B)*(E*A)*(D*C))"),
    .INIT(64'ha3330333a0000000))
    al_c6f13ae6 (
    .a(al_cc14f446),
    .b(al_473186ca),
    .c(al_2e8ff7ab),
    .d(al_54f03dbf[1]),
    .e(al_4f1a9685),
    .f(al_735aa681),
    .o(al_f7483e6d));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    al_5c42f8ed (
    .a(al_6cdf2816),
    .b(al_9907ae47),
    .c(al_aac09418[0]),
    .o(al_73eb08b7[0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_1f72baf2 (
    .a(al_2e8ff7ab),
    .b(al_77df94be),
    .c(al_e06bfe23),
    .d(al_535d21bf),
    .o(al_6cdf2816));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_8e558ad (
    .a(al_6cdf2816),
    .b(al_aac09418[0]),
    .c(al_aac09418[1]),
    .o(al_3370be13));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_84d1cf1e (
    .a(al_3370be13),
    .b(al_aac09418[2]),
    .c(al_aac09418[3]),
    .d(al_aac09418[4]),
    .o(al_c1d58f9c));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_6d4edc76 (
    .a(al_aac09418[5]),
    .b(al_aac09418[6]),
    .c(al_aac09418[7]),
    .d(al_aac09418[8]),
    .o(al_7557c0dc));
  AL_MAP_LUT5 #(
    .EQN("(~C*(E@(D*B*A)))"),
    .INIT(32'h070f0800))
    al_dbc1757a (
    .a(al_c1d58f9c),
    .b(al_7557c0dc),
    .c(al_9907ae47),
    .d(al_aac09418[9]),
    .e(al_aac09418[10]),
    .o(al_73eb08b7[10]));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*~A)))"),
    .INIT(16'h2310))
    al_c633f3fe (
    .a(al_6cdf2816),
    .b(al_9907ae47),
    .c(al_aac09418[0]),
    .d(al_aac09418[1]),
    .o(al_73eb08b7[1]));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_9f4527a2 (
    .a(al_3370be13),
    .b(al_9907ae47),
    .c(al_aac09418[2]),
    .o(al_73eb08b7[2]));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_b00be93d (
    .a(al_3370be13),
    .b(al_9907ae47),
    .c(al_aac09418[2]),
    .d(al_aac09418[3]),
    .o(al_73eb08b7[3]));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_5581fcce (
    .a(al_3370be13),
    .b(al_9907ae47),
    .c(al_aac09418[2]),
    .d(al_aac09418[3]),
    .e(al_aac09418[4]),
    .o(al_73eb08b7[4]));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    al_1f9564b1 (
    .a(al_c1d58f9c),
    .b(al_9907ae47),
    .c(al_aac09418[5]),
    .o(al_73eb08b7[5]));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_990b1cb0 (
    .a(al_c1d58f9c),
    .b(al_9907ae47),
    .c(al_aac09418[5]),
    .d(al_aac09418[6]),
    .o(al_73eb08b7[6]));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    al_13585585 (
    .a(al_c1d58f9c),
    .b(al_9907ae47),
    .c(al_aac09418[5]),
    .d(al_aac09418[6]),
    .e(al_aac09418[7]),
    .o(al_73eb08b7[7]));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F@(E*D*C*A)))"),
    .INIT(64'h1333333320000000))
    al_a356449e (
    .a(al_c1d58f9c),
    .b(al_9907ae47),
    .c(al_aac09418[5]),
    .d(al_aac09418[6]),
    .e(al_aac09418[7]),
    .f(al_aac09418[8]),
    .o(al_73eb08b7[8]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D@(B*A)))"),
    .INIT(16'h0708))
    al_9b415cba (
    .a(al_c1d58f9c),
    .b(al_7557c0dc),
    .c(al_9907ae47),
    .d(al_aac09418[9]),
    .o(al_73eb08b7[9]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_58959fda (
    .a(al_14016c23[3]),
    .b(al_aac09418[3]),
    .o(al_467061b3));
  AL_MAP_LUT6 #(
    .EQN("(B*A*~(F@D)*~(E@C))"),
    .INIT(64'h8000080000800008))
    al_7cd165fc (
    .a(al_be034ab5),
    .b(al_99f08586),
    .c(al_14016c23[5]),
    .d(al_14016c23[7]),
    .e(al_aac09418[5]),
    .f(al_aac09418[7]),
    .o(al_f205e138));
  AL_MAP_LUT6 #(
    .EQN("(~B*(F*~((A*~(E*~D)))*~(C)+F*(A*~(E*~D))*~(C)+~(F)*(A*~(E*~D))*C+F*(A*~(E*~D))*C))"),
    .INIT(64'h2303232320002020))
    al_a743e54a (
    .a(al_f205e138),
    .b(al_9907ae47),
    .c(al_77df94be),
    .d(al_14016c23[4]),
    .e(al_aac09418[4]),
    .f(al_994b00c4),
    .o(al_18337cf7));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_f3b11326 (
    .a(al_14016c23[6]),
    .b(al_aac09418[6]),
    .o(al_b42812f4));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(~E*B)*~(~D*A))"),
    .INIT(64'hf05030100f050301))
    al_47bef9db (
    .a(al_14016c23[0]),
    .b(al_14016c23[9]),
    .c(al_14016c23[10]),
    .d(al_aac09418[0]),
    .e(al_aac09418[9]),
    .f(al_aac09418[10]),
    .o(al_99f08586));
  AL_MAP_LUT6 #(
    .EQN("(~(~F*C)*~(E@B)*~(D*~A))"),
    .INIT(64'h88cc2233080c0203))
    al_324b8c3c (
    .a(al_14016c23[1]),
    .b(al_14016c23[2]),
    .c(al_14016c23[4]),
    .d(al_aac09418[1]),
    .e(al_aac09418[2]),
    .f(al_aac09418[4]),
    .o(al_bba5a10a));
  AL_MAP_LUT6 #(
    .EQN("(~(F@C)*~(~E*B)*~(D*~A))"),
    .INIT(64'ha0f020300a0f0203))
    al_50df2f07 (
    .a(al_14016c23[0]),
    .b(al_14016c23[1]),
    .c(al_14016c23[8]),
    .d(al_aac09418[0]),
    .e(al_aac09418[1]),
    .f(al_aac09418[8]),
    .o(al_70b7c327));
  AL_MAP_LUT6 #(
    .EQN("(~D*~C*B*A*~(F*~E))"),
    .INIT(64'h0008000000080008))
    al_38e9160f (
    .a(al_bba5a10a),
    .b(al_70b7c327),
    .c(al_467061b3),
    .d(al_b42812f4),
    .e(al_14016c23[9]),
    .f(al_aac09418[9]),
    .o(al_be034ab5));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_228e07f5 (
    .a(al_d86c9f70),
    .b(al_d1451a79),
    .o(al_618737cb));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    al_c24c6167 (
    .a(al_b242ee60[3]),
    .b(al_b242ee60[4]),
    .c(al_b242ee60[5]),
    .d(al_b242ee60[6]),
    .e(al_b242ee60[7]),
    .o(al_890eb5a1));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    al_80f611a1 (
    .a(al_d632949b),
    .b(al_2e8ff7ab),
    .c(al_54f03dbf[1]),
    .d(al_a783ebfd),
    .o(al_4290d1b8));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*B*A)"),
    .INIT(32'h00000080))
    al_673a6bb6 (
    .a(al_890eb5a1),
    .b(al_4290d1b8),
    .c(al_b242ee60[0]),
    .d(al_b242ee60[1]),
    .e(al_b242ee60[2]),
    .o(al_f0947bb5));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    al_99c5a530 (
    .a(al_890eb5a1),
    .b(al_b242ee60[0]),
    .c(al_b242ee60[1]),
    .d(al_b242ee60[2]),
    .o(al_d86c9f70));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_cfa649f1 (
    .a(al_d86c9f70),
    .b(al_4290d1b8),
    .o(al_8996909b));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(~D*~A))"),
    .INIT(16'h3f2a))
    al_853e8b6d (
    .a(al_473186ca),
    .b(al_d1ddae16),
    .c(al_e06bfe23),
    .d(al_fe00f314),
    .o(al_e1409b5e));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(D*~C*~B))"),
    .INIT(16'habaa))
    al_ad449554 (
    .a(al_473186ca),
    .b(al_9907ae47),
    .c(al_2ff03e70),
    .d(al_db3c8a2c),
    .o(al_a0088870));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_434ed8d7 (
    .a(al_603ec03),
    .b(al_7701781b),
    .o(al_473186ca));
  AL_MAP_LUT6 #(
    .EQN("(F*~E*~D*~A*~(C*B))"),
    .INIT(64'h0000001500000000))
    al_849afb9a (
    .a(al_9907ae47),
    .b(al_77df94be),
    .c(al_2ff03e70),
    .d(al_51ab8bb8),
    .e(al_1ed21a96),
    .f(al_2c7a1247),
    .o(al_2787c2b9));
  AL_MAP_LUT5 #(
    .EQN("~(~B*~(A*~(~E*D*~C)))"),
    .INIT(32'heeeeecee))
    al_7cd3f3cf (
    .a(al_2787c2b9),
    .b(al_473186ca),
    .c(al_d632949b),
    .d(al_994b00c4),
    .e(al_cca5b6a5),
    .o(al_4cf5bca0));
  AL_MAP_LUT6 #(
    .EQN("((F*~D*~C*~B)*~(E)*~(A)+(F*~D*~C*~B)*E*~(A)+~((F*~D*~C*~B))*E*A+(F*~D*~C*~B)*E*A)"),
    .INIT(64'haaab0001aaaa0000))
    al_d774b774 (
    .a(al_c5bc3747),
    .b(al_9907ae47),
    .c(al_535d21bf),
    .d(al_51ab8bb8),
    .e(al_fe00f314),
    .f(al_2c7a1247),
    .o(al_a396e89f));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_fe314073 (
    .a(al_2e8ff7ab),
    .b(al_54f03dbf[0]),
    .o(al_d1451a79));
  AL_MAP_LUT6 #(
    .EQN("~((~F*~B)*~((A*~(E*D)))*~(C)+(~F*~B)*(A*~(E*D))*~(C)+~((~F*~B))*(A*~(E*D))*C+(~F*~B)*(A*~(E*D))*C)"),
    .INIT(64'hff5f5f5ffc5c5c5c))
    al_63199624 (
    .a(al_890eb5a1),
    .b(al_473186ca),
    .c(al_d1451a79),
    .d(al_b242ee60[1]),
    .e(al_b242ee60[2]),
    .f(al_cca5b6a5),
    .o(al_63101725));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_ad61bd71 (
    .a(al_6ec43dd2),
    .b(al_1ff7640d),
    .o(al_949a133d));
  AL_MAP_LUT6 #(
    .EQN("((D*~B)*~((A*~(~F*~E)))*~(C)+(D*~B)*(A*~(~F*~E))*~(C)+~((D*~B))*(A*~(~F*~E))*C+(D*~B)*(A*~(~F*~E))*C)"),
    .INIT(64'ha3a0a3a0a3a00300))
    al_794d97db (
    .a(al_cc14f446),
    .b(al_9907ae47),
    .c(al_4f1a9685),
    .d(al_823fecd4),
    .e(al_8399b753),
    .f(al_88c53423),
    .o(al_27161c58));
  AL_DFF_X al_7c7c44cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0afd253[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(al_ff9a7266),
    .q(al_14016c23[0]));
  AL_DFF_X al_f1a94863 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0afd253[9]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(al_ff9a7266),
    .q(al_14016c23[9]));
  AL_DFF_X al_d0d0fd29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0afd253[10]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(al_ff9a7266),
    .q(al_14016c23[10]));
  AL_DFF_X al_a0cd6e4e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0afd253[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(al_ff9a7266),
    .q(al_14016c23[1]));
  AL_DFF_X al_d94145cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0afd253[2]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(al_ff9a7266),
    .q(al_14016c23[2]));
  AL_DFF_X al_ee326c34 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0afd253[3]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(al_ff9a7266),
    .q(al_14016c23[3]));
  AL_DFF_X al_6a162578 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0afd253[4]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(al_ff9a7266),
    .q(al_14016c23[4]));
  AL_DFF_X al_76fb5176 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0afd253[5]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(al_ff9a7266),
    .q(al_14016c23[5]));
  AL_DFF_X al_53c45e63 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0afd253[6]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(al_ff9a7266),
    .q(al_14016c23[6]));
  AL_DFF_X al_7f61f185 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0afd253[7]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(al_ff9a7266),
    .q(al_14016c23[7]));
  AL_DFF_X al_a6d6d77f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0afd253[8]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(al_ff9a7266),
    .q(al_14016c23[8]));
  AL_DFF_X al_d5116ac3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_73eb08b7[0]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_aac09418[0]));
  AL_DFF_X al_74e951f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_73eb08b7[9]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_aac09418[9]));
  AL_DFF_X al_f98d189c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_73eb08b7[10]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_aac09418[10]));
  AL_DFF_X al_4ca88e55 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_73eb08b7[1]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_aac09418[1]));
  AL_DFF_X al_5e4110f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_73eb08b7[2]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_aac09418[2]));
  AL_DFF_X al_2f5953a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_73eb08b7[3]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_aac09418[3]));
  AL_DFF_X al_dc853c99 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_73eb08b7[4]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_aac09418[4]));
  AL_DFF_X al_60716a49 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_73eb08b7[5]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_aac09418[5]));
  AL_DFF_X al_ea98976b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_73eb08b7[6]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_aac09418[6]));
  AL_DFF_X al_b0d7a40a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_73eb08b7[7]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_aac09418[7]));
  AL_DFF_X al_37f44914 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_73eb08b7[8]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_aac09418[8]));
  AL_DFF_X al_ec4685ea (
    .ar(al_ff9a7266),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_92477e6d[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cbc62139[0]));
  AL_DFF_X al_ca382286 (
    .ar(al_ff9a7266),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_92477e6d[9]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cbc62139[9]));
  AL_DFF_X al_ef5d1e05 (
    .ar(al_ff9a7266),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_92477e6d[10]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cbc62139[10]));
  AL_DFF_X al_6e5e9922 (
    .ar(al_ff9a7266),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_92477e6d[11]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cbc62139[11]));
  AL_DFF_X al_eaea2d3d (
    .ar(al_ff9a7266),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_92477e6d[12]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cbc62139[12]));
  AL_DFF_X al_82a11d37 (
    .ar(al_ff9a7266),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_92477e6d[13]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cbc62139[13]));
  AL_DFF_X al_4e9b0acc (
    .ar(al_ff9a7266),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_92477e6d[14]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cbc62139[14]));
  AL_DFF_X al_63594b3a (
    .ar(al_ff9a7266),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_92477e6d[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cbc62139[1]));
  AL_DFF_X al_23f155c7 (
    .ar(al_ff9a7266),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_92477e6d[2]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cbc62139[2]));
  AL_DFF_X al_6a4bcfe5 (
    .ar(al_ff9a7266),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_92477e6d[3]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cbc62139[3]));
  AL_DFF_X al_ff0f59fa (
    .ar(al_ff9a7266),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_92477e6d[4]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cbc62139[4]));
  AL_DFF_X al_b99fc69e (
    .ar(al_ff9a7266),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_92477e6d[5]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cbc62139[5]));
  AL_DFF_X al_6e9c07bb (
    .ar(al_ff9a7266),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_92477e6d[6]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cbc62139[6]));
  AL_DFF_X al_38474746 (
    .ar(al_ff9a7266),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_92477e6d[7]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cbc62139[7]));
  AL_DFF_X al_a7bcd582 (
    .ar(al_ff9a7266),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_92477e6d[8]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cbc62139[8]));
  AL_DFF_X al_282dbaa5 (
    .ar(al_ff9a7266),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_cbc62139[0]),
    .en(al_e7a9a14d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1f0d50be[0]));
  AL_DFF_X al_bd9c67ca (
    .ar(al_ff9a7266),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_cbc62139[9]),
    .en(al_e7a9a14d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1f0d50be[9]));
  AL_DFF_X al_2b024a13 (
    .ar(al_ff9a7266),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_cbc62139[10]),
    .en(al_e7a9a14d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1f0d50be[10]));
  AL_DFF_X al_ed070381 (
    .ar(al_ff9a7266),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_cbc62139[11]),
    .en(al_e7a9a14d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1f0d50be[11]));
  AL_DFF_X al_470eead5 (
    .ar(al_ff9a7266),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_cbc62139[12]),
    .en(al_e7a9a14d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1f0d50be[12]));
  AL_DFF_X al_7f90849f (
    .ar(al_ff9a7266),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_cbc62139[13]),
    .en(al_e7a9a14d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1f0d50be[13]));
  AL_DFF_X al_6f3a0d7 (
    .ar(al_ff9a7266),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_cbc62139[1]),
    .en(al_e7a9a14d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1f0d50be[1]));
  AL_DFF_X al_41aebefb (
    .ar(al_ff9a7266),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_cbc62139[2]),
    .en(al_e7a9a14d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1f0d50be[2]));
  AL_DFF_X al_4e8dcb15 (
    .ar(al_ff9a7266),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_cbc62139[3]),
    .en(al_e7a9a14d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1f0d50be[3]));
  AL_DFF_X al_d2459928 (
    .ar(al_ff9a7266),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_cbc62139[4]),
    .en(al_e7a9a14d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1f0d50be[4]));
  AL_DFF_X al_45b80aa0 (
    .ar(al_ff9a7266),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_cbc62139[5]),
    .en(al_e7a9a14d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1f0d50be[5]));
  AL_DFF_X al_90dd451a (
    .ar(al_ff9a7266),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_cbc62139[6]),
    .en(al_e7a9a14d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1f0d50be[6]));
  AL_DFF_X al_cd78758 (
    .ar(al_ff9a7266),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_cbc62139[7]),
    .en(al_e7a9a14d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1f0d50be[7]));
  AL_DFF_X al_e2036afd (
    .ar(al_ff9a7266),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_cbc62139[8]),
    .en(al_e7a9a14d),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1f0d50be[8]));
  AL_DFF_X al_1b495dda (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_87b441ee),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_d6a2be89[0]));
  AL_DFF_X al_f8901edb (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_59c37d06),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_d6a2be89[1]));
  AL_DFF_X al_a04c53c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f7f8cae),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_1feb4c09));
  AL_DFF_X al_ec9d500d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_90c946f9),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_54d691ed));
  AL_MAP_LUT5 #(
    .EQN("~(~C*~(D*~(E)*~((B*A))+D*E*~((B*A))+~(D)*E*(B*A)+D*E*(B*A)))"),
    .INIT(32'hfff8f7f0))
    al_76ede0db (
    .a(al_bbb4d320),
    .b(rx_clk_en),
    .c(al_ff9a7266),
    .d(al_54d691ed),
    .e(al_a0f12bef[2]),
    .o(al_90c946f9));
  AL_DFF_X al_67b07fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_34784d5d),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_f16920e0));
  AL_DFF_X al_99e6e826 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_68634068),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ff67665e));
  AL_MAP_LUT5 #(
    .EQN("(~C*(D*~(E)*~((B*A))+D*E*~((B*A))+~(D)*E*(B*A)+D*E*(B*A)))"),
    .INIT(32'h0f080700))
    al_2490cdb9 (
    .a(al_473186ca),
    .b(rx_clk_en),
    .c(al_ff9a7266),
    .d(al_ff67665e),
    .e(al_a0f12bef[5]),
    .o(al_68634068));
  AL_DFF_X al_a161f34c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e202820f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d632949b));
  AL_MAP_LUT5 #(
    .EQN("(~C*(D*~(E)*~((B*A))+D*E*~((B*A))+~(D)*E*(B*A)+D*E*(B*A)))"),
    .INIT(32'h0f080700))
    al_1833a7ac (
    .a(al_473186ca),
    .b(rx_clk_en),
    .c(al_ff9a7266),
    .d(al_d632949b),
    .e(al_a0f12bef[6]),
    .o(al_e202820f));
  AL_DFF_X al_2315c608 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_c702b161),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cc4e6731));
  AL_MAP_LUT5 #(
    .EQN("(~C*(D*~(E)*~((B*A))+D*E*~((B*A))+~(D)*E*(B*A)+D*E*(B*A)))"),
    .INIT(32'h0f080700))
    al_8d036bbc (
    .a(al_473186ca),
    .b(rx_clk_en),
    .c(al_ff9a7266),
    .d(al_cc4e6731),
    .e(al_a0f12bef[7]),
    .o(al_c702b161));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    al_dc4e2f6c (
    .a(al_4b9a6e34),
    .b(al_f4c47e2b[3]),
    .c(al_4c524efc[3]),
    .d(al_93bf05b4[3]),
    .o(al_34784d5d));
  AL_DFF_X al_22f890a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_46f5ce71),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_7bce675b));
  AL_DFF_X al_4f31b55d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_7bce675b),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_f9cac200));
  AL_DFF_X al_4f23830b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_8867ef3c[2]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_a7a7af9e));
  AL_DFF_X al_6bb0e19e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_a7a7af9e),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_c2569e9f));
  AL_DFF_X al_70ddf8f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_89fbca82),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_d0a10128));
  AL_DFF_X al_e0cf31ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_628888c[3]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_3da78c22));
  AL_DFF_X al_da8c7197 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_3da78c22),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_db0897ce));
  AL_DFF_X al_f6c44eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_29f8870a),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_e06bfe23));
  AL_DFF_X al_31262525 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_89eb3505),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_77df94be));
  AL_DFF_X al_45f4b890 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1a86743a),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_d5b2f5c4));
  AL_DFF_X al_1839851a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b3eb9d64),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_2ff03e70));
  AL_DFF_X al_a327e535 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_77be5888),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_6627cbad));
  AL_DFF_X al_314476ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_289fe017),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_d1ddae16));
  AL_DFF_X al_7a0f4a21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_7f375c7a),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_9907ae47));
  AL_DFF_X al_1fd0276a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_abc7ca1f),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_535d21bf));
  AL_DFF_X al_13ee25a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_db547825),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_2e8ff7ab));
  AL_DFF_X al_eca9de50 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_6bfa7885),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_7701781b));
  AL_DFF_X al_ac073428 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_8f82c138),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_614db0a6));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_6b758b67 (
    .a(al_4b9a6e34),
    .b(al_f4c47e2b[3]),
    .c(al_4c524efc[3]),
    .d(al_93bf05b4[3]),
    .o(al_2f3f17d));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~(C*~B*~A))"),
    .INIT(32'h00ef0000))
    al_a92e1327 (
    .a(al_2f3f17d),
    .b(al_8867ef3c[2]),
    .c(al_628888c[3]),
    .d(al_6627cbad),
    .e(al_535d21bf),
    .o(al_77be5888));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_da685628 (
    .a(al_7bce675b),
    .b(al_f9cac200),
    .o(al_b3eb9d64));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    al_d10e0719 (
    .a(al_d57700f8[3]),
    .b(al_d5e21796[3]),
    .c(al_8867ef3c[2]),
    .d(al_628888c[3]),
    .o(al_c1e4e3b));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    al_74cfcf9f (
    .a(al_c1e4e3b),
    .b(al_f6dc28d8[3]),
    .c(al_5d5249da[3]),
    .d(al_ba4af77d[3]),
    .o(al_4b9a6e34));
  AL_MAP_LUT6 #(
    .EQN("(~F*~A*~(~E*~(D*~C*~B)))"),
    .INIT(64'h0000000055550100))
    al_47c16cbe (
    .a(al_49bc5cf4),
    .b(al_c2569e9f),
    .c(al_3da78c22),
    .d(al_db0897ce),
    .e(al_6627cbad),
    .f(al_9907ae47),
    .o(al_67caff7a));
  AL_MAP_LUT6 #(
    .EQN("(C*~B*~(A*(~(D)*~(E)*~(F)+D*E*F)))"),
    .INIT(64'h1030303030303010))
    al_e5586377 (
    .a(al_4b9a6e34),
    .b(al_49bc5cf4),
    .c(al_3da78c22),
    .d(al_f4c47e2b[3]),
    .e(al_4c524efc[3]),
    .f(al_93bf05b4[3]),
    .o(al_5ae0e8ee));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~(D*~C*~A))"),
    .INIT(16'hcdcc))
    al_37582bf2 (
    .a(al_5ae0e8ee),
    .b(al_67caff7a),
    .c(al_a7a7af9e),
    .d(al_c2569e9f),
    .o(al_7f375c7a));
  AL_MAP_LUT5 #(
    .EQN("(B*~(~(E*~D)*~(~C*A)))"),
    .INIT(32'h08cc0808))
    al_8e2b2d97 (
    .a(al_316af0f0),
    .b(al_a7a7af9e),
    .c(al_c2569e9f),
    .d(al_603ec03),
    .e(al_7701781b),
    .o(al_6bfa7885));
  AL_MAP_LUT6 #(
    .EQN("(~F*A*~(~E*~(C*~(~D*B))))"),
    .INIT(64'h00000000aaaaa020))
    al_918c0624 (
    .a(al_a7a7af9e),
    .b(al_c2569e9f),
    .c(al_603ec03),
    .d(al_7701781b),
    .e(al_d5b2f5c4),
    .f(al_54f03dbf[5]),
    .o(al_1a86743a));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT(16'h88a0))
    al_1479574d (
    .a(al_a7a7af9e),
    .b(al_d5b2f5c4),
    .c(al_614db0a6),
    .d(al_54f03dbf[5]),
    .o(al_8f82c138));
  AL_MAP_LUT5 #(
    .EQN("(~D*A*~(~C*~(E*B)))"),
    .INIT(32'h00a800a0))
    al_36fdbc68 (
    .a(al_a7a7af9e),
    .b(al_614db0a6),
    .c(al_2e8ff7ab),
    .d(al_54f03dbf[1]),
    .e(al_54f03dbf[5]),
    .o(al_db547825));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_308b5b13 (
    .a(al_a7a7af9e),
    .b(al_8867ef3c[2]),
    .o(al_289fe017));
  AL_MAP_LUT5 #(
    .EQN("(~E*A*~(~C*~(D*B)))"),
    .INIT(32'h0000a8a0))
    al_47029a9d (
    .a(al_a7a7af9e),
    .b(al_2e8ff7ab),
    .c(al_77df94be),
    .d(al_54f03dbf[1]),
    .e(al_2ff03e70),
    .o(al_89eb3505));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*~A))"),
    .INIT(8'hf4))
    al_a326183a (
    .a(al_d1ddae16),
    .b(al_e06bfe23),
    .c(al_2ff03e70),
    .o(al_29f8870a));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_bbe73f5 (
    .a(al_a7a7af9e),
    .b(al_3da78c22),
    .o(al_e8517c4));
  AL_MAP_LUT6 #(
    .EQN("(~D*~C*~B*A*~(~F*~E))"),
    .INIT(64'h0002000200020000))
    al_f4f9ef89 (
    .a(al_e8517c4),
    .b(al_49bc5cf4),
    .c(al_f16920e0),
    .d(al_6ecd5054),
    .e(al_e06bfe23),
    .f(al_535d21bf),
    .o(al_abc7ca1f));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~A*~(~E*~D*~C*~B))"),
    .INIT(64'hffffffffaaaaaaab))
    al_6ac46427 (
    .a(al_9907ae47),
    .b(al_d5b2f5c4),
    .c(al_614db0a6),
    .d(al_2e8ff7ab),
    .e(al_e06bfe23),
    .f(al_54f03dbf[5]),
    .o(al_71b48cc2[0]));
  AL_MAP_LUT6 #(
    .EQN("(F*~A*~(~E*~D*~C*~B))"),
    .INIT(64'h5555555400000000))
    al_543f4750 (
    .a(al_9907ae47),
    .b(al_d5b2f5c4),
    .c(al_614db0a6),
    .d(al_2e8ff7ab),
    .e(al_e06bfe23),
    .f(al_54f03dbf[0]),
    .o(al_71b48cc2[1]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_9c1780c5 (
    .a(al_9907ae47),
    .b(al_54f03dbf[1]),
    .o(al_516522f9[0]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_e637ff22 (
    .a(al_9907ae47),
    .b(al_54f03dbf[2]),
    .o(al_516522f9[1]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_4c6b9740 (
    .a(al_9907ae47),
    .b(al_54f03dbf[3]),
    .o(al_516522f9[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_368b9d64 (
    .a(al_9907ae47),
    .b(al_54f03dbf[4]),
    .o(al_516522f9[3]));
  AL_DFF_X al_b7a123bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_71b48cc2[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(al_ff9a7266),
    .q(al_54f03dbf[0]));
  AL_DFF_X al_9b59c0a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_71b48cc2[1]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_54f03dbf[1]));
  AL_DFF_X al_e7e41b85 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_516522f9[0]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_54f03dbf[2]));
  AL_DFF_X al_4b0bf56f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_516522f9[1]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_54f03dbf[3]));
  AL_DFF_X al_4bb7e3f3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_516522f9[2]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_54f03dbf[4]));
  AL_DFF_X al_e3561075 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_516522f9[3]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_54f03dbf[5]));
  AL_DFF_X al_deeffd93 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_43bf9cc4),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_status_vld));
  AL_DFF_X al_3b2a8f5a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_921d9eff),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_603ec03));
  AL_DFF_X al_c35e88c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_321e78bf),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49bc5cf4));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(~D*~(E)*~((B*A))+~D*E*~((B*A))+~(~D)*E*(B*A)+~D*E*(B*A)))"),
    .INIT(32'h07000f08))
    al_4e3513c (
    .a(al_473186ca),
    .b(rx_clk_en),
    .c(al_ff9a7266),
    .d(al_49bc5cf4),
    .e(al_25215c55[1]),
    .o(al_321e78bf));
  AL_DFF_X al_6d42a679 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_6c890ee8),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_43bf9cc4));
  AL_DFF_X al_efe7003c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_a87a1c23),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_d280e871));
  AL_DFF_X al_b0a4c438 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_3119a20d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_531e5772));
  AL_MAP_LUT5 #(
    .EQN("(~C*(D*~(E)*~((B*A))+D*E*~((B*A))+~(D)*E*(B*A)+D*E*(B*A)))"),
    .INIT(32'h0f080700))
    al_5da6ee97 (
    .a(al_473186ca),
    .b(rx_clk_en),
    .c(al_ff9a7266),
    .d(al_531e5772),
    .e(al_a0f12bef[3]),
    .o(al_3119a20d));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_1c0afab6 (
    .a(al_d280e871),
    .b(al_cd9c4b15),
    .o(al_f7f8cae));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_caa7289c (
    .a(al_d280e871),
    .b(al_a14eea73),
    .o(al_3e7ed8af));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_776f7d7e (
    .a(al_5772dfd3),
    .b(al_e4bdca8a),
    .o(al_b1b61f7c[0]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_1173f73e (
    .a(al_5772dfd3),
    .b(al_e4bdca8a),
    .o(al_b1b61f7c[1]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    al_61fa61fe (
    .a(al_a7a7af9e),
    .b(al_3da78c22),
    .c(al_4b3fffb5[1]),
    .d(al_4b3fffb5[3]),
    .o(al_da5fd7db));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_632220af (
    .a(al_da5fd7db),
    .b(al_4b3fffb5[4]),
    .c(al_4b3fffb5[6]),
    .d(al_4b3fffb5[7]),
    .o(al_80344ab4));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    al_309aa20b (
    .a(al_80344ab4),
    .b(al_4b3fffb5[0]),
    .c(al_4b3fffb5[2]),
    .d(al_4b3fffb5[5]),
    .o(al_921d9eff));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*C*B*A)"),
    .INIT(64'h0000000000000080))
    al_49bbf960 (
    .a(al_e8517c4),
    .b(al_4b3fffb5[1]),
    .c(al_4b3fffb5[3]),
    .d(al_4b3fffb5[4]),
    .e(al_4b3fffb5[6]),
    .f(al_4b3fffb5[7]),
    .o(al_749e1728));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    al_820d44bb (
    .a(al_749e1728),
    .b(al_4b3fffb5[0]),
    .c(al_4b3fffb5[2]),
    .d(al_4b3fffb5[5]),
    .o(al_6baf9e53));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    al_e2053c (
    .a(al_e8c5f626[0]),
    .b(al_e8c5f626[2]),
    .c(al_e8c5f626[4]),
    .d(al_e8c5f626[6]),
    .e(al_e8c5f626[7]),
    .o(al_7bee3de4));
  AL_MAP_LUT6 #(
    .EQN("(~F*~(~E*~D*~C*~B*A))"),
    .INIT(64'h00000000fffffffd))
    al_9ce063c1 (
    .a(al_7bee3de4),
    .b(al_d0a10128),
    .c(al_e8c5f626[1]),
    .d(al_e8c5f626[3]),
    .e(al_e8c5f626[5]),
    .f(al_9e8909aa),
    .o(al_8d11b694));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_6210d2b5 (
    .a(al_8d11b694),
    .b(al_7bce675b),
    .o(al_3252df70));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_172766e8 (
    .a(al_ad22e376),
    .b(al_4596a396),
    .o(al_59a83809));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~(~B*~(C*A)))"),
    .INIT(32'h000000ec))
    al_9a4852b6 (
    .a(al_59a83809),
    .b(al_d280e871),
    .c(al_cac2565f),
    .d(al_cd9c4b15),
    .e(al_a14eea73),
    .o(al_a87a1c23));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    al_2fa3367b (
    .a(al_59a83809),
    .b(al_d280e871),
    .c(al_cac2565f),
    .o(al_6281ecee));
  AL_DFF_X al_b27fbca0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_cd9c4b15),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_c5802d0a[0]));
  AL_DFF_X al_ed8c264c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1f0d50be[4]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_c5802d0a[9]));
  AL_DFF_X al_e630ab06 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1f0d50be[5]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_c5802d0a[10]));
  AL_DFF_X al_e69ed9b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1f0d50be[6]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_c5802d0a[11]));
  AL_DFF_X al_fb35ff7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1f0d50be[7]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_c5802d0a[12]));
  AL_DFF_X al_d56664e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1f0d50be[8]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_c5802d0a[13]));
  AL_DFF_X al_4a16db11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1f0d50be[9]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_c5802d0a[14]));
  AL_DFF_X al_8b470712 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1f0d50be[10]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_c5802d0a[15]));
  AL_DFF_X al_dbca1a9d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1f0d50be[11]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_c5802d0a[16]));
  AL_DFF_X al_69788c51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1f0d50be[12]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_c5802d0a[17]));
  AL_DFF_X al_d5a91f1d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1f0d50be[13]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_c5802d0a[18]));
  AL_DFF_X al_d16cc316 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_a14eea73),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_c5802d0a[1]));
  AL_DFF_X al_f13c369f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_8e811a01),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_c5802d0a[19]));
  AL_DFF_X al_85c1c6ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_dc6fb7d9),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_c5802d0a[20]));
  AL_DFF_X al_b2a6d110 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_391ec013),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_c5802d0a[21]));
  AL_DFF_X al_f850d904 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_32839ce1),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_c5802d0a[23]));
  AL_DFF_X al_b9b8940e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b1b61f7c[1]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_c5802d0a[24]));
  AL_DFF_X al_b55f70b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b1b61f7c[0]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_c5802d0a[2]));
  AL_DFF_X al_7ce2f40b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_9f0e53e2[5]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_c5802d0a[3]));
  AL_DFF_X al_d5c516ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ed990b15),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_c5802d0a[4]));
  AL_DFF_X al_4211f31f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1f0d50be[0]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_c5802d0a[5]));
  AL_DFF_X al_670c0085 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1f0d50be[1]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_c5802d0a[6]));
  AL_DFF_X al_9f77adcb (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1f0d50be[2]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_c5802d0a[7]));
  AL_DFF_X al_10f3f751 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1f0d50be[3]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_c5802d0a[8]));
  AL_DFF_X al_11693e9c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_fa90a029[0]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_e8c5f626[0]));
  AL_DFF_X al_41058574 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_fa90a029[1]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_e8c5f626[1]));
  AL_DFF_X al_bea0dfa3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_fa90a029[2]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_e8c5f626[2]));
  AL_DFF_X al_96ca5ab2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_fa90a029[3]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_e8c5f626[3]));
  AL_DFF_X al_8b926098 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_fa90a029[4]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_e8c5f626[4]));
  AL_DFF_X al_e243cfa1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_fa90a029[5]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_e8c5f626[5]));
  AL_DFF_X al_648c8e20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_fa90a029[6]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_e8c5f626[6]));
  AL_DFF_X al_923d20ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_fa90a029[7]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_e8c5f626[7]));
  AL_DFF_X al_364014d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ba4af77d[3]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_4b3fffb5[0]));
  AL_DFF_X al_5bd03593 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_93bf05b4[3]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_4b3fffb5[1]));
  AL_DFF_X al_14f0914a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_4c524efc[3]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_4b3fffb5[2]));
  AL_DFF_X al_5f12d685 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f4c47e2b[3]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_4b3fffb5[3]));
  AL_DFF_X al_18477828 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5d5249da[3]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_4b3fffb5[4]));
  AL_DFF_X al_441b00d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f6dc28d8[3]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_4b3fffb5[5]));
  AL_DFF_X al_d735eed0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_d5e21796[3]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_4b3fffb5[6]));
  AL_DFF_X al_5a13c9f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_d57700f8[3]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_4b3fffb5[7]));
  AL_DFF_X al_a0e1de1f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_4b3fffb5[0]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_b242ee60[0]));
  AL_DFF_X al_f1c0b0e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_4b3fffb5[1]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_b242ee60[1]));
  AL_DFF_X al_7ee0d1df (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_4b3fffb5[2]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_b242ee60[2]));
  AL_DFF_X al_188f0d62 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_4b3fffb5[3]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_b242ee60[3]));
  AL_DFF_X al_6e6d04f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_4b3fffb5[4]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_b242ee60[4]));
  AL_DFF_X al_faaca9ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_4b3fffb5[5]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_b242ee60[5]));
  AL_DFF_X al_2834fadc (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_4b3fffb5[6]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_b242ee60[6]));
  AL_DFF_X al_6ca7503f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_4b3fffb5[7]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_b242ee60[7]));
  AL_DFF_X al_7180eafe (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b242ee60[0]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_12d2a17a[0]));
  AL_DFF_X al_d54eedbb (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b242ee60[1]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_12d2a17a[1]));
  AL_DFF_X al_73bf3bee (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b242ee60[2]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_12d2a17a[2]));
  AL_DFF_X al_74371668 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b242ee60[3]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_12d2a17a[3]));
  AL_DFF_X al_b9328f65 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b242ee60[4]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_12d2a17a[4]));
  AL_DFF_X al_5955628e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b242ee60[5]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_12d2a17a[5]));
  AL_DFF_X al_79d20d73 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b242ee60[6]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_12d2a17a[6]));
  AL_DFF_X al_e6f90e56 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_b242ee60[7]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_12d2a17a[7]));
  AL_DFF_X al_e1095791 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_12d2a17a[0]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_5160c8c2[0]));
  AL_DFF_X al_fd4f17d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_12d2a17a[1]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_5160c8c2[1]));
  AL_DFF_X al_aee85b3c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_12d2a17a[2]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_5160c8c2[2]));
  AL_DFF_X al_507114da (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_12d2a17a[3]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_5160c8c2[3]));
  AL_DFF_X al_67357f5a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_12d2a17a[4]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_5160c8c2[4]));
  AL_DFF_X al_e80e8480 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_12d2a17a[5]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_5160c8c2[5]));
  AL_DFF_X al_d7551ee5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_12d2a17a[6]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_5160c8c2[6]));
  AL_DFF_X al_a7f0057b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_12d2a17a[7]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_5160c8c2[7]));
  AL_DFF_X al_2fa377f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_c5802d0a[0]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_status_vector[0]));
  AL_DFF_X al_d5b96e06 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_c5802d0a[9]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_status_vector[9]));
  AL_DFF_X al_af9f446 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_c5802d0a[10]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_status_vector[10]));
  AL_DFF_X al_651ffa98 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_c5802d0a[11]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_status_vector[11]));
  AL_DFF_X al_df9c40cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_c5802d0a[12]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_status_vector[12]));
  AL_DFF_X al_62cbdab6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_c5802d0a[13]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_status_vector[13]));
  AL_DFF_X al_af40b71 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_c5802d0a[14]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_status_vector[14]));
  AL_DFF_X al_ff642eb2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_c5802d0a[15]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_status_vector[15]));
  AL_DFF_X al_11c6f619 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_c5802d0a[16]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_status_vector[16]));
  AL_DFF_X al_58df1fd5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_c5802d0a[17]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_status_vector[17]));
  AL_DFF_X al_2d5f2ea9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_c5802d0a[18]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_status_vector[18]));
  AL_DFF_X al_21f27d75 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_c5802d0a[1]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_status_vector[1]));
  AL_DFF_X al_2b0aea47 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_c5802d0a[19]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_status_vector[21]));
  AL_DFF_X al_ce0f2315 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_c5802d0a[20]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_status_vector[19]));
  AL_DFF_X al_ba0ed298 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_c5802d0a[21]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_status_vector[22]));
  AL_DFF_X al_9e0f29e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_c5802d0a[23]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_status_vector[20]));
  AL_DFF_X al_ac774633 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_c5802d0a[24]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_status_vector[25]));
  AL_DFF_X al_b8d4022d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_c5802d0a[2]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_status_vector[26]));
  AL_DFF_X al_36f5528b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_c5802d0a[3]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_status_vector[2]));
  AL_DFF_X al_8e1e439b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_c5802d0a[4]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_status_vector[3]));
  AL_DFF_X al_9fa723a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_c5802d0a[5]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_status_vector[5]));
  AL_DFF_X al_429e0317 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_c5802d0a[6]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_status_vector[6]));
  AL_DFF_X al_fcb54c8b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_c5802d0a[7]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_status_vector[7]));
  AL_DFF_X al_409284d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_c5802d0a[8]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_status_vector[8]));
  AL_DFF_0 al_82d24448 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e8c5f626[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ba4af77d[0]));
  AL_DFF_0 al_490a6dc7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ba4af77d[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ba4af77d[1]));
  AL_DFF_0 al_be8f3415 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ba4af77d[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ba4af77d[2]));
  AL_DFF_0 al_28ab72ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ba4af77d[2]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ba4af77d[3]));
  AL_DFF_0 al_2b108e65 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e8c5f626[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_93bf05b4[0]));
  AL_DFF_0 al_f047df1a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_93bf05b4[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_93bf05b4[1]));
  AL_DFF_0 al_a897a45f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_93bf05b4[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_93bf05b4[2]));
  AL_DFF_0 al_e7d35e9e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_93bf05b4[2]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_93bf05b4[3]));
  AL_DFF_0 al_9f80cec0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e8c5f626[2]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c524efc[0]));
  AL_DFF_0 al_fe9e922a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_4c524efc[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c524efc[1]));
  AL_DFF_0 al_9db09235 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_4c524efc[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c524efc[2]));
  AL_DFF_0 al_b7d88b91 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_4c524efc[2]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c524efc[3]));
  AL_DFF_0 al_a87f8afe (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e8c5f626[3]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f4c47e2b[0]));
  AL_DFF_0 al_dd0e6243 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f4c47e2b[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f4c47e2b[1]));
  AL_DFF_0 al_47e3702d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f4c47e2b[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f4c47e2b[2]));
  AL_DFF_0 al_62fad1f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f4c47e2b[2]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f4c47e2b[3]));
  AL_DFF_0 al_ec2fe39f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e8c5f626[4]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5d5249da[0]));
  AL_DFF_0 al_36d86ddb (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5d5249da[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5d5249da[1]));
  AL_DFF_0 al_4457e5b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5d5249da[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5d5249da[2]));
  AL_DFF_0 al_eb6e6159 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_5d5249da[2]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5d5249da[3]));
  AL_DFF_0 al_f45bd9a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e8c5f626[5]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f6dc28d8[0]));
  AL_DFF_0 al_22d81463 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f6dc28d8[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f6dc28d8[1]));
  AL_DFF_0 al_f2d5653e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f6dc28d8[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f6dc28d8[2]));
  AL_DFF_0 al_2687c550 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f6dc28d8[2]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f6dc28d8[3]));
  AL_DFF_0 al_aef5aabc (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e8c5f626[6]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d5e21796[0]));
  AL_DFF_0 al_f312af84 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_d5e21796[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d5e21796[1]));
  AL_DFF_0 al_b46ca986 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_d5e21796[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d5e21796[2]));
  AL_DFF_0 al_efddb838 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_d5e21796[2]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d5e21796[3]));
  AL_DFF_0 al_cabbf2bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_e8c5f626[7]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d57700f8[0]));
  AL_DFF_0 al_f4cf992f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_d57700f8[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d57700f8[1]));
  AL_DFF_0 al_db440685 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_d57700f8[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d57700f8[2]));
  AL_DFF_0 al_d572d894 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_d57700f8[2]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d57700f8[3]));
  AL_DFF_X al_a2a8bbff (
    .ar(1'b0),
    .as(al_1e2edecf),
    .clk(rx_mac_clk),
    .d(1'b0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e18a88b8));
  AL_DFF_X al_6f236533 (
    .ar(1'b0),
    .as(al_1e2edecf),
    .clk(rx_mac_clk),
    .d(al_e18a88b8),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fcf500fb));
  AL_DFF_X al_80374e42 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_fcf500fb),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7f87fb2e));
  AL_DFF_X al_6eefe3b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_fc3fb77f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ff9a7266));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_537c02db (
    .a(al_fcf500fb),
    .b(al_7f87fb2e),
    .o(al_fc3fb77f));
  AL_DFF_X al_55ac0271 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_72f5321b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(speed_100));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    al_6a02fd2c (
    .a(al_25215c55[1]),
    .o(al_61aea43e));
  AL_DFF_X al_ec87a88 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_61aea43e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6ea32e9c));
  AL_DFF_X al_42e988dc (
    .ar(1'b0),
    .as(al_6d2cc211),
    .clk(tx_mac_clk),
    .d(1'b0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3f3dfbd));
  AL_DFF_X al_4bf1b3b0 (
    .ar(1'b0),
    .as(al_6d2cc211),
    .clk(tx_mac_clk),
    .d(al_d3f3dfbd),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2a91cf37));
  AL_DFF_X al_343bc1fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2a91cf37),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f13f5376));
  AL_DFF_X al_552d4cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9fe1548f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6b4499fc));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_1c9ced9 (
    .a(al_2a91cf37),
    .b(al_f13f5376),
    .o(al_9fe1548f));
  AL_MAP_LUT4 #(
    .EQN("((D*~B)*~(C)*~(A)+(D*~B)*C*~(A)+~((D*~B))*C*A+(D*~B)*C*A)"),
    .INIT(16'hb1a0))
    al_f5710c5a (
    .a(tx_clk_en),
    .b(al_6b4499fc),
    .c(al_ae5f998b[0]),
    .d(al_ae5f998b[1]),
    .o(al_e1759dc[0]));
  AL_MAP_LUT4 #(
    .EQN("((D*~B)*~(C)*~(A)+(D*~B)*C*~(A)+~((D*~B))*C*A+(D*~B)*C*A)"),
    .INIT(16'hb1a0))
    al_c8792b39 (
    .a(tx_clk_en),
    .b(al_6b4499fc),
    .c(al_ae5f998b[10]),
    .d(al_ae5f998b[11]),
    .o(al_e1759dc[10]));
  AL_MAP_LUT4 #(
    .EQN("((D*~B)*~(C)*~(A)+(D*~B)*C*~(A)+~((D*~B))*C*A+(D*~B)*C*A)"),
    .INIT(16'hb1a0))
    al_8ec8c0a (
    .a(tx_clk_en),
    .b(al_6b4499fc),
    .c(al_ae5f998b[11]),
    .d(al_ae5f998b[12]),
    .o(al_e1759dc[11]));
  AL_MAP_LUT4 #(
    .EQN("((D*~B)*~(C)*~(A)+(D*~B)*C*~(A)+~((D*~B))*C*A+(D*~B)*C*A)"),
    .INIT(16'hb1a0))
    al_a9b6604c (
    .a(tx_clk_en),
    .b(al_6b4499fc),
    .c(al_ae5f998b[12]),
    .d(al_ae5f998b[13]),
    .o(al_e1759dc[12]));
  AL_MAP_LUT4 #(
    .EQN("((D*~B)*~(C)*~(A)+(D*~B)*C*~(A)+~((D*~B))*C*A+(D*~B)*C*A)"),
    .INIT(16'hb1a0))
    al_dbe7a94b (
    .a(tx_clk_en),
    .b(al_6b4499fc),
    .c(al_ae5f998b[13]),
    .d(al_ae5f998b[14]),
    .o(al_e1759dc[13]));
  AL_MAP_LUT4 #(
    .EQN("((D*~B)*~(C)*~(A)+(D*~B)*C*~(A)+~((D*~B))*C*A+(D*~B)*C*A)"),
    .INIT(16'hb1a0))
    al_387c06db (
    .a(tx_clk_en),
    .b(al_6b4499fc),
    .c(al_ae5f998b[1]),
    .d(al_ae5f998b[2]),
    .o(al_e1759dc[1]));
  AL_MAP_LUT4 #(
    .EQN("((D*~B)*~(C)*~(A)+(D*~B)*C*~(A)+~((D*~B))*C*A+(D*~B)*C*A)"),
    .INIT(16'hb1a0))
    al_567dee6 (
    .a(tx_clk_en),
    .b(al_6b4499fc),
    .c(al_ae5f998b[2]),
    .d(al_ae5f998b[3]),
    .o(al_e1759dc[2]));
  AL_MAP_LUT4 #(
    .EQN("((D*~B)*~(C)*~(A)+(D*~B)*C*~(A)+~((D*~B))*C*A+(D*~B)*C*A)"),
    .INIT(16'hb1a0))
    al_c03f5970 (
    .a(tx_clk_en),
    .b(al_6b4499fc),
    .c(al_ae5f998b[3]),
    .d(al_ae5f998b[4]),
    .o(al_e1759dc[3]));
  AL_MAP_LUT4 #(
    .EQN("((D*~B)*~(C)*~(A)+(D*~B)*C*~(A)+~((D*~B))*C*A+(D*~B)*C*A)"),
    .INIT(16'hb1a0))
    al_a81e1d04 (
    .a(tx_clk_en),
    .b(al_6b4499fc),
    .c(al_ae5f998b[4]),
    .d(al_ae5f998b[5]),
    .o(al_e1759dc[4]));
  AL_MAP_LUT4 #(
    .EQN("((D*~B)*~(C)*~(A)+(D*~B)*C*~(A)+~((D*~B))*C*A+(D*~B)*C*A)"),
    .INIT(16'hb1a0))
    al_4efb6f27 (
    .a(tx_clk_en),
    .b(al_6b4499fc),
    .c(al_ae5f998b[5]),
    .d(al_ae5f998b[6]),
    .o(al_e1759dc[5]));
  AL_MAP_LUT4 #(
    .EQN("((D*~B)*~(C)*~(A)+(D*~B)*C*~(A)+~((D*~B))*C*A+(D*~B)*C*A)"),
    .INIT(16'hb1a0))
    al_51970e96 (
    .a(tx_clk_en),
    .b(al_6b4499fc),
    .c(al_ae5f998b[6]),
    .d(al_ae5f998b[7]),
    .o(al_e1759dc[6]));
  AL_MAP_LUT4 #(
    .EQN("((D*~B)*~(C)*~(A)+(D*~B)*C*~(A)+~((D*~B))*C*A+(D*~B)*C*A)"),
    .INIT(16'hb1a0))
    al_74b9fe3b (
    .a(tx_clk_en),
    .b(al_6b4499fc),
    .c(al_ae5f998b[7]),
    .d(al_ae5f998b[8]),
    .o(al_e1759dc[7]));
  AL_MAP_LUT4 #(
    .EQN("((D*~B)*~(C)*~(A)+(D*~B)*C*~(A)+~((D*~B))*C*A+(D*~B)*C*A)"),
    .INIT(16'hb1a0))
    al_4bd2820f (
    .a(tx_clk_en),
    .b(al_6b4499fc),
    .c(al_ae5f998b[8]),
    .d(al_ae5f998b[9]),
    .o(al_e1759dc[8]));
  AL_MAP_LUT4 #(
    .EQN("((D*~B)*~(C)*~(A)+(D*~B)*C*~(A)+~((D*~B))*C*A+(D*~B)*C*A)"),
    .INIT(16'hb1a0))
    al_176f504c (
    .a(tx_clk_en),
    .b(al_6b4499fc),
    .c(al_ae5f998b[9]),
    .d(al_ae5f998b[10]),
    .o(al_e1759dc[9]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_e6df14e5 (
    .a(al_ae5f998b[13]),
    .b(al_ae5f998b[14]),
    .o(al_dc745a17));
  AL_DFF_X al_a0d3b26a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_dc745a17),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_ae5f998b[0]));
  AL_DFF_X al_ee9240ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e1759dc[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ae5f998b[9]));
  AL_DFF_X al_7e871877 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e1759dc[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ae5f998b[10]));
  AL_DFF_X al_c8fb12f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e1759dc[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ae5f998b[11]));
  AL_DFF_X al_e9d559ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e1759dc[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ae5f998b[12]));
  AL_DFF_X al_de380fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e1759dc[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ae5f998b[13]));
  AL_DFF_X al_b8f0e9ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e1759dc[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ae5f998b[14]));
  AL_DFF_X al_e41223f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e1759dc[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ae5f998b[1]));
  AL_DFF_X al_b0f1ad03 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e1759dc[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ae5f998b[2]));
  AL_DFF_X al_eef3b243 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e1759dc[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ae5f998b[3]));
  AL_DFF_X al_55fa39b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e1759dc[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ae5f998b[4]));
  AL_DFF_X al_f2828325 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e1759dc[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ae5f998b[5]));
  AL_DFF_X al_b99eb840 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e1759dc[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ae5f998b[6]));
  AL_DFF_X al_e1e00dd8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e1759dc[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ae5f998b[7]));
  AL_DFF_X al_2c2b9e9e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e1759dc[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ae5f998b[8]));
  AL_DFF_X al_653c0943 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ae5f998b[14]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_6c9db937[0]));
  AL_DFF_X al_88a7e11d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_6c9db937[8]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_6c9db937[9]));
  AL_DFF_X al_3417e8c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_6c9db937[0]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_6c9db937[1]));
  AL_DFF_X al_5eac4751 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_6c9db937[1]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_6c9db937[2]));
  AL_DFF_X al_925e636e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_6c9db937[2]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_6c9db937[3]));
  AL_DFF_X al_61d8a91c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_6c9db937[3]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_6c9db937[4]));
  AL_DFF_X al_98dd875f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_6c9db937[4]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_6c9db937[5]));
  AL_DFF_X al_68c66282 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_6c9db937[5]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_6c9db937[6]));
  AL_DFF_X al_bac6a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_6c9db937[6]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_6c9db937[7]));
  AL_DFF_X al_c16c8f4f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_6c9db937[7]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_6c9db937[8]));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(~D*~C*B))"),
    .INIT(16'h555d))
    al_16e67e73 (
    .a(al_ed1f021e[0]),
    .b(al_e702d1c[0]),
    .c(al_e702d1c[1]),
    .d(al_e702d1c[2]),
    .o(al_3a9d8027[0]));
  AL_MAP_LUT5 #(
    .EQN("(~(~E*~D*C)*~(B@A))"),
    .INIT(32'h99999909))
    al_508b5ec (
    .a(al_ed1f021e[0]),
    .b(al_ed1f021e[1]),
    .c(al_e702d1c[0]),
    .d(al_e702d1c[1]),
    .e(al_e702d1c[2]),
    .o(al_3a9d8027[1]));
  AL_MAP_LUT6 #(
    .EQN("~(~(~F*~E*D)*~(C@(~B*~A)))"),
    .INIT(64'he1e1e1e1e1e1ffe1))
    al_246499ee (
    .a(al_ed1f021e[0]),
    .b(al_ed1f021e[1]),
    .c(al_ed1f021e[2]),
    .d(al_e702d1c[0]),
    .e(al_e702d1c[1]),
    .f(al_e702d1c[2]),
    .o(al_3a9d8027[2]));
  AL_MAP_LUT4 #(
    .EQN("~(D@(~C*~B*~A))"),
    .INIT(16'h01fe))
    al_1fa38748 (
    .a(al_ed1f021e[0]),
    .b(al_ed1f021e[1]),
    .c(al_ed1f021e[2]),
    .d(al_ed1f021e[3]),
    .o(al_3d691a71));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~D*~C*B))"),
    .INIT(16'h5551))
    al_bd9154f9 (
    .a(al_3d691a71),
    .b(al_e702d1c[0]),
    .c(al_e702d1c[1]),
    .d(al_e702d1c[2]),
    .o(al_3a9d8027[3]));
  AL_MAP_LUT5 #(
    .EQN("~(E*~(C)*~((~D*~B*~A))+E*C*~((~D*~B*~A))+~(E)*C*(~D*~B*~A)+E*C*(~D*~B*~A))"),
    .INIT(32'h0001ffef))
    al_38d5e436 (
    .a(al_ed1f021e[0]),
    .b(al_ed1f021e[1]),
    .c(al_ed1f021e[2]),
    .d(al_ed1f021e[3]),
    .e(al_e702d1c[0]),
    .o(al_c9a41ba));
  AL_MAP_LUT6 #(
    .EQN("(~E*(~(A)*~(C)*D*~((F*B))+~(A)*C*D*~((F*B))+~(A)*~(C)*~(D)*(F*B)+A*~(C)*~(D)*(F*B)+~(A)*C*~(D)*(F*B)+A*C*~(D)*(F*B)+~(A)*~(C)*D*(F*B)+A*~(C)*D*(F*B)+~(A)*C*D*(F*B)))"),
    .INIT(64'h00005dcc00005500))
    al_86547198 (
    .a(al_c9a41ba),
    .b(al_977227b4),
    .c(al_e702d1c[0]),
    .d(al_e702d1c[1]),
    .e(al_e702d1c[2]),
    .f(al_9b4eaefc[2]),
    .o(al_536d34[0]));
  AL_MAP_LUT6 #(
    .EQN("(~E*(~(A)*C*~(D)*~((F*B))+A*C*~(D)*~((F*B))+~(A)*~(C)*D*~((F*B))+A*~(C)*D*~((F*B))+~(A)*C*D*~((F*B))+~(A)*C*D*(F*B)))"),
    .INIT(64'h0000533000005ff0))
    al_621229cd (
    .a(al_eccfd98c),
    .b(al_977227b4),
    .c(al_e702d1c[0]),
    .d(al_e702d1c[1]),
    .e(al_e702d1c[2]),
    .f(al_9b4eaefc[2]),
    .o(al_536d34[1]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_37a2f086 (
    .a(al_ed1f021e[0]),
    .b(al_ed1f021e[1]),
    .c(al_ed1f021e[2]),
    .d(al_ed1f021e[3]),
    .o(al_eccfd98c));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E)"),
    .INIT(32'h000ca000))
    al_cd90c74c (
    .a(al_eccfd98c),
    .b(al_7cd73f8f),
    .c(al_e702d1c[0]),
    .d(al_e702d1c[1]),
    .e(al_e702d1c[2]),
    .o(al_536d34[2]));
  AL_DFF_X al_76403bf8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_3a9d8027[0]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_ed1f021e[0]));
  AL_DFF_X al_26be93f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_3a9d8027[1]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_ed1f021e[1]));
  AL_DFF_X al_4ec4e657 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_3a9d8027[2]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_ed1f021e[2]));
  AL_DFF_X al_2fc90547 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_3a9d8027[3]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_ed1f021e[3]));
  AL_DFF_X al_864e1fb1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_536d34[0]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_e702d1c[0]));
  AL_DFF_X al_de9aedd5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_536d34[1]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_e702d1c[1]));
  AL_DFF_X al_43028ed6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_536d34[2]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_e702d1c[2]));
  AL_DFF_X al_2e5c085 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2c5269c),
    .en(al_a162bb8e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_beea368e));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_40ed4686 (
    .a(tx_clk_en),
    .b(al_6b4499fc),
    .o(al_a162bb8e));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_d1fa6c25 (
    .a(al_2337d80f),
    .b(al_10fc4c0e),
    .c(al_edc29fee),
    .o(al_3c42ccfe));
  AL_MAP_LUT5 #(
    .EQN("(~E*~C*~(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))"),
    .INIT(32'h0000050c))
    al_673b1263 (
    .a(al_5ef35ad0),
    .b(al_3c42ccfe),
    .c(al_ea30f787),
    .d(al_b01f953d[0]),
    .e(al_b01f953d[1]),
    .o(al_ed15c12c[0]));
  AL_MAP_LUT6 #(
    .EQN("(A*~((~D*~C*B))*E*~(F)+A*(~D*~C*B)*E*~(F)+~(A)*(~D*~C*B)*~(E)*F+A*(~D*~C*B)*~(E)*F)"),
    .INIT(64'h0000000caaaa0000))
    al_d359a3e1 (
    .a(al_5ef35ad0),
    .b(al_2337d80f),
    .c(al_ea30f787),
    .d(al_cf085f09),
    .e(al_b01f953d[0]),
    .f(al_b01f953d[1]),
    .o(al_ed15c12c[1]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~A*~(~D*~B)))"),
    .INIT(16'ha0b0))
    al_cb38e35 (
    .a(al_beea368e),
    .b(al_715819dc[4]),
    .c(al_b01f953d[0]),
    .d(al_b01f953d[1]),
    .o(al_2c5269c));
  AL_MAP_LUT6 #(
    .EQN("(~((~B*~A))*~(C)*~(D)*~(E)*~(F)+(~B*~A)*~(C)*~(D)*~(E)*~(F)+~((~B*~A))*C*~(D)*~(E)*~(F)+(~B*~A)*C*~(D)*~(E)*~(F)+~((~B*~A))*~(C)*D*~(E)*~(F)+(~B*~A)*~(C)*D*~(E)*~(F)+~((~B*~A))*C*D*~(E)*~(F)+(~B*~A)*C*D*~(E)*~(F)+(~B*~A)*C*~(D)*E*~(F)+~((~B*~A))*~(C)*D*E*~(F)+~((~B*~A))*C*D*E*~(F)+(~B*~A)*C*D*E*~(F)+~((~B*~A))*~(C)*D*~(E)*F+(~B*~A)*~(C)*D*~(E)*F+~((~B*~A))*C*D*~(E)*F+(~B*~A)*C*D*~(E)*F+~((~B*~A))*~(C)*D*E*F+(~B*~A)*~(C)*D*E*F+~((~B*~A))*C*D*E*F+(~B*~A)*C*D*E*F)"),
    .INIT(64'hff00ff00fe10ffff))
    al_cad392d6 (
    .a(al_5ef35ad0),
    .b(al_ea30f787),
    .c(al_72a2cf60[0]),
    .d(al_715819dc[0]),
    .e(al_b01f953d[0]),
    .f(al_b01f953d[1]),
    .o(al_1f1bbfc9[0]));
  AL_MAP_LUT6 #(
    .EQN("(~((~B*~A))*~(C)*~(D)*~(E)*~(F)+(~B*~A)*~(C)*~(D)*~(E)*~(F)+~((~B*~A))*C*~(D)*~(E)*~(F)+(~B*~A)*C*~(D)*~(E)*~(F)+~((~B*~A))*~(C)*D*~(E)*~(F)+(~B*~A)*~(C)*D*~(E)*~(F)+~((~B*~A))*C*D*~(E)*~(F)+(~B*~A)*C*D*~(E)*~(F)+(~B*~A)*C*~(D)*E*~(F)+~((~B*~A))*~(C)*D*E*~(F)+~((~B*~A))*C*D*E*~(F)+(~B*~A)*C*D*E*~(F)+~((~B*~A))*~(C)*D*~(E)*F+(~B*~A)*~(C)*D*~(E)*F+~((~B*~A))*C*D*~(E)*F+(~B*~A)*C*D*~(E)*F+~((~B*~A))*~(C)*D*E*F+(~B*~A)*~(C)*D*E*F+~((~B*~A))*C*D*E*F+(~B*~A)*C*D*E*F)"),
    .INIT(64'hff00ff00fe10ffff))
    al_6c157c7b (
    .a(al_5ef35ad0),
    .b(al_ea30f787),
    .c(al_72a2cf60[10]),
    .d(al_715819dc[10]),
    .e(al_b01f953d[0]),
    .f(al_b01f953d[1]),
    .o(al_1f1bbfc9[10]));
  AL_MAP_LUT6 #(
    .EQN("(~((~B*~A))*~(C)*~(D)*~(E)*~(F)+(~B*~A)*~(C)*~(D)*~(E)*~(F)+~((~B*~A))*C*~(D)*~(E)*~(F)+(~B*~A)*C*~(D)*~(E)*~(F)+~((~B*~A))*~(C)*D*~(E)*~(F)+(~B*~A)*~(C)*D*~(E)*~(F)+~((~B*~A))*C*D*~(E)*~(F)+(~B*~A)*C*D*~(E)*~(F)+(~B*~A)*C*~(D)*E*~(F)+~((~B*~A))*~(C)*D*E*~(F)+~((~B*~A))*C*D*E*~(F)+(~B*~A)*C*D*E*~(F)+~((~B*~A))*~(C)*D*~(E)*F+(~B*~A)*~(C)*D*~(E)*F+~((~B*~A))*C*D*~(E)*F+(~B*~A)*C*D*~(E)*F+~((~B*~A))*~(C)*D*E*F+(~B*~A)*~(C)*D*E*F+~((~B*~A))*C*D*E*F+(~B*~A)*C*D*E*F)"),
    .INIT(64'hff00ff00fe10ffff))
    al_1f3b189c (
    .a(al_5ef35ad0),
    .b(al_ea30f787),
    .c(al_72a2cf60[11]),
    .d(al_715819dc[11]),
    .e(al_b01f953d[0]),
    .f(al_b01f953d[1]),
    .o(al_1f1bbfc9[11]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_95733d66 (
    .a(al_715819dc[0]),
    .b(al_715819dc[1]),
    .c(al_715819dc[2]),
    .d(al_715819dc[3]),
    .e(al_715819dc[4]),
    .f(al_715819dc[5]),
    .o(al_46fe62ca));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_f8fada65 (
    .a(al_715819dc[6]),
    .b(al_715819dc[7]),
    .c(al_715819dc[8]),
    .d(al_715819dc[9]),
    .o(al_c504b787));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    al_fe7a523c (
    .a(al_46fe62ca),
    .b(al_c504b787),
    .c(al_715819dc[10]),
    .d(al_715819dc[11]),
    .e(al_715819dc[12]),
    .o(al_5ef35ad0));
  AL_MAP_LUT6 #(
    .EQN("(~((~B*~A))*~(C)*~(D)*~(E)*~(F)+(~B*~A)*~(C)*~(D)*~(E)*~(F)+~((~B*~A))*C*~(D)*~(E)*~(F)+(~B*~A)*C*~(D)*~(E)*~(F)+~((~B*~A))*~(C)*D*~(E)*~(F)+(~B*~A)*~(C)*D*~(E)*~(F)+~((~B*~A))*C*D*~(E)*~(F)+(~B*~A)*C*D*~(E)*~(F)+(~B*~A)*C*~(D)*E*~(F)+~((~B*~A))*~(C)*D*E*~(F)+~((~B*~A))*C*D*E*~(F)+(~B*~A)*C*D*E*~(F)+~((~B*~A))*~(C)*D*~(E)*F+(~B*~A)*~(C)*D*~(E)*F+~((~B*~A))*C*D*~(E)*F+(~B*~A)*C*D*~(E)*F+~((~B*~A))*~(C)*D*E*F+(~B*~A)*~(C)*D*E*F+~((~B*~A))*C*D*E*F+(~B*~A)*C*D*E*F)"),
    .INIT(64'hff00ff00fe10ffff))
    al_b03e19ed (
    .a(al_5ef35ad0),
    .b(al_ea30f787),
    .c(al_72a2cf60[12]),
    .d(al_715819dc[12]),
    .e(al_b01f953d[0]),
    .f(al_b01f953d[1]),
    .o(al_1f1bbfc9[12]));
  AL_MAP_LUT6 #(
    .EQN("(~((~B*~A))*~(C)*~(D)*~(E)*~(F)+(~B*~A)*~(C)*~(D)*~(E)*~(F)+~((~B*~A))*C*~(D)*~(E)*~(F)+(~B*~A)*C*~(D)*~(E)*~(F)+~((~B*~A))*~(C)*D*~(E)*~(F)+(~B*~A)*~(C)*D*~(E)*~(F)+~((~B*~A))*C*D*~(E)*~(F)+(~B*~A)*C*D*~(E)*~(F)+(~B*~A)*C*~(D)*E*~(F)+~((~B*~A))*~(C)*D*E*~(F)+~((~B*~A))*C*D*E*~(F)+(~B*~A)*C*D*E*~(F)+~((~B*~A))*~(C)*D*~(E)*F+(~B*~A)*~(C)*D*~(E)*F+~((~B*~A))*C*D*~(E)*F+(~B*~A)*C*D*~(E)*F+~((~B*~A))*~(C)*D*E*F+(~B*~A)*~(C)*D*E*F+~((~B*~A))*C*D*E*F+(~B*~A)*C*D*E*F)"),
    .INIT(64'hff00ff00fe10ffff))
    al_33d5c5a4 (
    .a(al_5ef35ad0),
    .b(al_ea30f787),
    .c(al_72a2cf60[1]),
    .d(al_715819dc[1]),
    .e(al_b01f953d[0]),
    .f(al_b01f953d[1]),
    .o(al_1f1bbfc9[1]));
  AL_MAP_LUT6 #(
    .EQN("(~((~B*~A))*~(C)*~(D)*~(E)*~(F)+(~B*~A)*~(C)*~(D)*~(E)*~(F)+~((~B*~A))*C*~(D)*~(E)*~(F)+(~B*~A)*C*~(D)*~(E)*~(F)+~((~B*~A))*~(C)*D*~(E)*~(F)+(~B*~A)*~(C)*D*~(E)*~(F)+~((~B*~A))*C*D*~(E)*~(F)+(~B*~A)*C*D*~(E)*~(F)+(~B*~A)*C*~(D)*E*~(F)+~((~B*~A))*~(C)*D*E*~(F)+~((~B*~A))*C*D*E*~(F)+(~B*~A)*C*D*E*~(F)+~((~B*~A))*~(C)*D*~(E)*F+(~B*~A)*~(C)*D*~(E)*F+~((~B*~A))*C*D*~(E)*F+(~B*~A)*C*D*~(E)*F+~((~B*~A))*~(C)*D*E*F+(~B*~A)*~(C)*D*E*F+~((~B*~A))*C*D*E*F+(~B*~A)*C*D*E*F)"),
    .INIT(64'hff00ff00fe10ffff))
    al_58131b99 (
    .a(al_5ef35ad0),
    .b(al_ea30f787),
    .c(al_72a2cf60[2]),
    .d(al_715819dc[2]),
    .e(al_b01f953d[0]),
    .f(al_b01f953d[1]),
    .o(al_1f1bbfc9[2]));
  AL_MAP_LUT6 #(
    .EQN("(~((~B*~A))*~(C)*~(D)*~(E)*~(F)+(~B*~A)*~(C)*~(D)*~(E)*~(F)+~((~B*~A))*C*~(D)*~(E)*~(F)+(~B*~A)*C*~(D)*~(E)*~(F)+~((~B*~A))*~(C)*D*~(E)*~(F)+(~B*~A)*~(C)*D*~(E)*~(F)+~((~B*~A))*C*D*~(E)*~(F)+(~B*~A)*C*D*~(E)*~(F)+(~B*~A)*C*~(D)*E*~(F)+~((~B*~A))*~(C)*D*E*~(F)+~((~B*~A))*C*D*E*~(F)+(~B*~A)*C*D*E*~(F)+~((~B*~A))*~(C)*D*~(E)*F+(~B*~A)*~(C)*D*~(E)*F+~((~B*~A))*C*D*~(E)*F+(~B*~A)*C*D*~(E)*F+~((~B*~A))*~(C)*D*E*F+(~B*~A)*~(C)*D*E*F+~((~B*~A))*C*D*E*F+(~B*~A)*C*D*E*F)"),
    .INIT(64'hff00ff00fe10ffff))
    al_8e35f97c (
    .a(al_5ef35ad0),
    .b(al_ea30f787),
    .c(al_72a2cf60[3]),
    .d(al_715819dc[3]),
    .e(al_b01f953d[0]),
    .f(al_b01f953d[1]),
    .o(al_1f1bbfc9[3]));
  AL_MAP_LUT6 #(
    .EQN("(~((~B*~A))*~(C)*~(D)*~(E)*~(F)+(~B*~A)*~(C)*~(D)*~(E)*~(F)+~((~B*~A))*C*~(D)*~(E)*~(F)+(~B*~A)*C*~(D)*~(E)*~(F)+~((~B*~A))*~(C)*D*~(E)*~(F)+(~B*~A)*~(C)*D*~(E)*~(F)+~((~B*~A))*C*D*~(E)*~(F)+(~B*~A)*C*D*~(E)*~(F)+(~B*~A)*C*~(D)*E*~(F)+~((~B*~A))*~(C)*D*E*~(F)+~((~B*~A))*C*D*E*~(F)+(~B*~A)*C*D*E*~(F)+~((~B*~A))*~(C)*D*~(E)*F+(~B*~A)*~(C)*D*~(E)*F+~((~B*~A))*C*D*~(E)*F+(~B*~A)*C*D*~(E)*F+~((~B*~A))*~(C)*D*E*F+(~B*~A)*~(C)*D*E*F+~((~B*~A))*C*D*E*F+(~B*~A)*C*D*E*F)"),
    .INIT(64'hff00ff00fe10ffff))
    al_26fe2456 (
    .a(al_5ef35ad0),
    .b(al_ea30f787),
    .c(al_72a2cf60[4]),
    .d(al_715819dc[4]),
    .e(al_b01f953d[0]),
    .f(al_b01f953d[1]),
    .o(al_1f1bbfc9[4]));
  AL_MAP_LUT6 #(
    .EQN("(~((~B*~A))*~(C)*~(D)*~(E)*~(F)+(~B*~A)*~(C)*~(D)*~(E)*~(F)+~((~B*~A))*C*~(D)*~(E)*~(F)+(~B*~A)*C*~(D)*~(E)*~(F)+~((~B*~A))*~(C)*D*~(E)*~(F)+(~B*~A)*~(C)*D*~(E)*~(F)+~((~B*~A))*C*D*~(E)*~(F)+(~B*~A)*C*D*~(E)*~(F)+(~B*~A)*C*~(D)*E*~(F)+~((~B*~A))*~(C)*D*E*~(F)+~((~B*~A))*C*D*E*~(F)+(~B*~A)*C*D*E*~(F)+~((~B*~A))*~(C)*D*~(E)*F+(~B*~A)*~(C)*D*~(E)*F+~((~B*~A))*C*D*~(E)*F+(~B*~A)*C*D*~(E)*F+~((~B*~A))*~(C)*D*E*F+(~B*~A)*~(C)*D*E*F+~((~B*~A))*C*D*E*F+(~B*~A)*C*D*E*F)"),
    .INIT(64'hff00ff00fe10ffff))
    al_b611d1bd (
    .a(al_5ef35ad0),
    .b(al_ea30f787),
    .c(al_72a2cf60[5]),
    .d(al_715819dc[5]),
    .e(al_b01f953d[0]),
    .f(al_b01f953d[1]),
    .o(al_1f1bbfc9[5]));
  AL_MAP_LUT6 #(
    .EQN("(~((~B*~A))*~(C)*~(D)*~(E)*~(F)+(~B*~A)*~(C)*~(D)*~(E)*~(F)+~((~B*~A))*C*~(D)*~(E)*~(F)+(~B*~A)*C*~(D)*~(E)*~(F)+~((~B*~A))*~(C)*D*~(E)*~(F)+(~B*~A)*~(C)*D*~(E)*~(F)+~((~B*~A))*C*D*~(E)*~(F)+(~B*~A)*C*D*~(E)*~(F)+(~B*~A)*C*~(D)*E*~(F)+~((~B*~A))*~(C)*D*E*~(F)+~((~B*~A))*C*D*E*~(F)+(~B*~A)*C*D*E*~(F)+~((~B*~A))*~(C)*D*~(E)*F+(~B*~A)*~(C)*D*~(E)*F+~((~B*~A))*C*D*~(E)*F+(~B*~A)*C*D*~(E)*F+~((~B*~A))*~(C)*D*E*F+(~B*~A)*~(C)*D*E*F+~((~B*~A))*C*D*E*F+(~B*~A)*C*D*E*F)"),
    .INIT(64'hff00ff00fe10ffff))
    al_4106cbf5 (
    .a(al_5ef35ad0),
    .b(al_ea30f787),
    .c(al_72a2cf60[6]),
    .d(al_715819dc[6]),
    .e(al_b01f953d[0]),
    .f(al_b01f953d[1]),
    .o(al_1f1bbfc9[6]));
  AL_MAP_LUT6 #(
    .EQN("(~((~B*~A))*~(C)*~(D)*~(E)*~(F)+(~B*~A)*~(C)*~(D)*~(E)*~(F)+~((~B*~A))*C*~(D)*~(E)*~(F)+(~B*~A)*C*~(D)*~(E)*~(F)+~((~B*~A))*~(C)*D*~(E)*~(F)+(~B*~A)*~(C)*D*~(E)*~(F)+~((~B*~A))*C*D*~(E)*~(F)+(~B*~A)*C*D*~(E)*~(F)+(~B*~A)*C*~(D)*E*~(F)+~((~B*~A))*~(C)*D*E*~(F)+~((~B*~A))*C*D*E*~(F)+(~B*~A)*C*D*E*~(F)+~((~B*~A))*~(C)*D*~(E)*F+(~B*~A)*~(C)*D*~(E)*F+~((~B*~A))*C*D*~(E)*F+(~B*~A)*C*D*~(E)*F+~((~B*~A))*~(C)*D*E*F+(~B*~A)*~(C)*D*E*F+~((~B*~A))*C*D*E*F+(~B*~A)*C*D*E*F)"),
    .INIT(64'hff00ff00fe10ffff))
    al_e5964cbf (
    .a(al_5ef35ad0),
    .b(al_ea30f787),
    .c(al_72a2cf60[7]),
    .d(al_715819dc[7]),
    .e(al_b01f953d[0]),
    .f(al_b01f953d[1]),
    .o(al_1f1bbfc9[7]));
  AL_MAP_LUT6 #(
    .EQN("(~((~B*~A))*~(C)*~(D)*~(E)*~(F)+(~B*~A)*~(C)*~(D)*~(E)*~(F)+~((~B*~A))*C*~(D)*~(E)*~(F)+(~B*~A)*C*~(D)*~(E)*~(F)+~((~B*~A))*~(C)*D*~(E)*~(F)+(~B*~A)*~(C)*D*~(E)*~(F)+~((~B*~A))*C*D*~(E)*~(F)+(~B*~A)*C*D*~(E)*~(F)+(~B*~A)*C*~(D)*E*~(F)+~((~B*~A))*~(C)*D*E*~(F)+~((~B*~A))*C*D*E*~(F)+(~B*~A)*C*D*E*~(F)+~((~B*~A))*~(C)*D*~(E)*F+(~B*~A)*~(C)*D*~(E)*F+~((~B*~A))*C*D*~(E)*F+(~B*~A)*C*D*~(E)*F+~((~B*~A))*~(C)*D*E*F+(~B*~A)*~(C)*D*E*F+~((~B*~A))*C*D*E*F+(~B*~A)*C*D*E*F)"),
    .INIT(64'hff00ff00fe10ffff))
    al_ad94922c (
    .a(al_5ef35ad0),
    .b(al_ea30f787),
    .c(al_72a2cf60[8]),
    .d(al_715819dc[8]),
    .e(al_b01f953d[0]),
    .f(al_b01f953d[1]),
    .o(al_1f1bbfc9[8]));
  AL_MAP_LUT6 #(
    .EQN("(~((~B*~A))*~(C)*~(D)*~(E)*~(F)+(~B*~A)*~(C)*~(D)*~(E)*~(F)+~((~B*~A))*C*~(D)*~(E)*~(F)+(~B*~A)*C*~(D)*~(E)*~(F)+~((~B*~A))*~(C)*D*~(E)*~(F)+(~B*~A)*~(C)*D*~(E)*~(F)+~((~B*~A))*C*D*~(E)*~(F)+(~B*~A)*C*D*~(E)*~(F)+(~B*~A)*C*~(D)*E*~(F)+~((~B*~A))*~(C)*D*E*~(F)+~((~B*~A))*C*D*E*~(F)+(~B*~A)*C*D*E*~(F)+~((~B*~A))*~(C)*D*~(E)*F+(~B*~A)*~(C)*D*~(E)*F+~((~B*~A))*C*D*~(E)*F+(~B*~A)*C*D*~(E)*F+~((~B*~A))*~(C)*D*E*F+(~B*~A)*~(C)*D*E*F+~((~B*~A))*C*D*E*F+(~B*~A)*C*D*E*F)"),
    .INIT(64'hff00ff00fe10ffff))
    al_d6271c13 (
    .a(al_5ef35ad0),
    .b(al_ea30f787),
    .c(al_72a2cf60[9]),
    .d(al_715819dc[9]),
    .e(al_b01f953d[0]),
    .f(al_b01f953d[1]),
    .o(al_1f1bbfc9[9]));
  AL_DFF_X al_39fdb056 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1f1bbfc9[0]),
    .en(al_a162bb8e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_715819dc[0]));
  AL_DFF_X al_d3f27480 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1f1bbfc9[9]),
    .en(al_a162bb8e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_715819dc[9]));
  AL_DFF_X al_54c0610d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1f1bbfc9[10]),
    .en(al_a162bb8e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_715819dc[10]));
  AL_DFF_X al_543ba014 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1f1bbfc9[11]),
    .en(al_a162bb8e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_715819dc[11]));
  AL_DFF_X al_93fd36e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1f1bbfc9[12]),
    .en(al_a162bb8e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_715819dc[12]));
  AL_DFF_X al_314d4832 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1f1bbfc9[1]),
    .en(al_a162bb8e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_715819dc[1]));
  AL_DFF_X al_4ec412c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1f1bbfc9[2]),
    .en(al_a162bb8e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_715819dc[2]));
  AL_DFF_X al_a95c96df (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1f1bbfc9[3]),
    .en(al_a162bb8e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_715819dc[3]));
  AL_DFF_X al_70d8f890 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1f1bbfc9[4]),
    .en(al_a162bb8e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_715819dc[4]));
  AL_DFF_X al_3a21f74a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1f1bbfc9[5]),
    .en(al_a162bb8e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_715819dc[5]));
  AL_DFF_X al_84e5c58a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1f1bbfc9[6]),
    .en(al_a162bb8e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_715819dc[6]));
  AL_DFF_X al_5dc14581 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1f1bbfc9[7]),
    .en(al_a162bb8e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_715819dc[7]));
  AL_DFF_X al_4e45259e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1f1bbfc9[8]),
    .en(al_a162bb8e),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_715819dc[8]));
  AL_DFF_X al_fd22e68d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ed15c12c[0]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_b01f953d[0]));
  AL_DFF_X al_65fd9e60 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ed15c12c[1]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_b01f953d[1]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_70a8eb70 (
    .a(1'b0),
    .o({al_eefcdfd,open_n10}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f2c3b06b (
    .a(al_715819dc[0]),
    .b(1'b1),
    .c(al_eefcdfd),
    .o({al_58846bb5,al_72a2cf60[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e71da01 (
    .a(al_715819dc[1]),
    .b(1'b0),
    .c(al_58846bb5),
    .o({al_6303158d,al_72a2cf60[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ee1be4ef (
    .a(al_715819dc[2]),
    .b(1'b0),
    .c(al_6303158d),
    .o({al_34d58259,al_72a2cf60[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_957049ca (
    .a(al_715819dc[3]),
    .b(1'b0),
    .c(al_34d58259),
    .o({al_69600a84,al_72a2cf60[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f8862321 (
    .a(al_715819dc[4]),
    .b(1'b0),
    .c(al_69600a84),
    .o({al_ebcb9742,al_72a2cf60[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c02bfe8e (
    .a(al_715819dc[5]),
    .b(1'b0),
    .c(al_ebcb9742),
    .o({al_7b06746d,al_72a2cf60[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e8284c3b (
    .a(al_715819dc[6]),
    .b(1'b0),
    .c(al_7b06746d),
    .o({al_bd268370,al_72a2cf60[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1a5f39ca (
    .a(al_715819dc[7]),
    .b(1'b0),
    .c(al_bd268370),
    .o({al_64206da8,al_72a2cf60[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f960a90d (
    .a(al_715819dc[8]),
    .b(1'b0),
    .c(al_64206da8),
    .o({al_922f69ff,al_72a2cf60[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4ddd0d7c (
    .a(al_715819dc[9]),
    .b(1'b0),
    .c(al_922f69ff),
    .o({al_baa25bac,al_72a2cf60[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_49fbabe1 (
    .a(al_715819dc[10]),
    .b(1'b0),
    .c(al_baa25bac),
    .o({al_22f4f2dd,al_72a2cf60[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f8a47967 (
    .a(al_715819dc[11]),
    .b(1'b0),
    .c(al_22f4f2dd),
    .o({al_7a3587c3,al_72a2cf60[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3f72ff06 (
    .a(al_715819dc[12]),
    .b(1'b0),
    .c(al_7a3587c3),
    .o({open_n11,al_72a2cf60[12]}));
  AL_DFF_X al_d8ab1b7f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_fadd6423),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_7ac4c27f));
  AL_DFF_X al_c8c45800 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(gmii_crs),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_977227b4));
  AL_DFF_X al_1234a145 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9b4eaefc[1]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_87969af9));
  AL_DFF_X al_e184f7a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9b4eaefc[2]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_10fc4c0e));
  AL_DFF_X al_3abf7331 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9b4eaefc[6]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_dd9e938b));
  AL_DFF_X al_cc372baa (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9b4eaefc[5]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_8cc75feb));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    al_7426b6e8 (
    .a(al_5f257019[2]),
    .o(al_e23c1f65[0]));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    al_8a2bb006 (
    .a(al_5f257019[3]),
    .o(al_e23c1f65[1]));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    al_fbd62836 (
    .a(al_5f257019[4]),
    .o(al_e23c1f65[2]));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    al_9f4b6d04 (
    .a(al_5f257019[5]),
    .o(al_e23c1f65[3]));
  AL_DFF_X al_53011a0d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_61aea43e),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_54081406));
  AL_DFF_X al_3c8b9f6b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_aa427d37),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_6b5283b3));
  AL_DFF_X al_fe622681 (
    .ar(al_6b4499fc),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_bc71f40f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4fb6999c));
  AL_MAP_LUT6 #(
    .EQN("(A*(B*~((~F*~E*~D))*~(C)+B*(~F*~E*~D)*~(C)+~(B)*(~F*~E*~D)*C+B*(~F*~E*~D)*C))"),
    .INIT(64'h08080808080808a8))
    al_ce366304 (
    .a(al_57798083),
    .b(al_1887f4c),
    .c(al_edc29fee),
    .d(al_e8bb9040[6]),
    .e(al_e8bb9040[7]),
    .f(al_e8bb9040[8]),
    .o(al_64ec9565));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*~B))"),
    .INIT(8'hba))
    al_88f7784d (
    .a(al_64ec9565),
    .b(tx_clk_en),
    .c(al_4fb6999c),
    .o(al_bc71f40f));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_45404119 (
    .a(al_e8bb9040[16]),
    .b(al_e8bb9040[17]),
    .c(al_e8bb9040[18]),
    .o(al_1887f4c));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*A)"),
    .INIT(64'h0000000000000002))
    al_4ed13ee7 (
    .a(tx_clk_en),
    .b(al_e8bb9040[3]),
    .c(al_e8bb9040[9]),
    .d(al_e8bb9040[10]),
    .e(al_e8bb9040[11]),
    .f(al_e8bb9040[12]),
    .o(al_ead880b8));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*A)"),
    .INIT(64'h0000000000000002))
    al_83882059 (
    .a(al_ead880b8),
    .b(al_e8bb9040[0]),
    .c(al_e8bb9040[1]),
    .d(al_e8bb9040[13]),
    .e(al_e8bb9040[14]),
    .f(al_e8bb9040[15]),
    .o(al_57798083));
  AL_DFF_X al_aefc4972 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f28fd6dc),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_c925873));
  AL_DFF_X al_13a6df02 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_af806095),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_a494216e));
  AL_DFF_X al_2d2f88c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ab89cd63),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_7fe117d0));
  AL_DFF_X al_aa7e42b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_3b1a77d7),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_e3f5d0d6));
  AL_DFF_X al_bb7b9aa3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4fe9a477),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_68ba43d4));
  AL_DFF_X al_c30ea28d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_df015ce6),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_12358921));
  AL_DFF_X al_cf6a05b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d277135),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_c2463579));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_a3bb5cb8 (
    .a(al_5411d218),
    .b(al_2a71f823),
    .c(al_8a6ca59e[0]),
    .o(al_a7d56e64[0]));
  AL_MAP_LUT3 #(
    .EQN("(C@(B*~A))"),
    .INIT(8'hb4))
    al_eaabfcb4 (
    .a(al_c78fe3c1),
    .b(al_2a71f823),
    .c(al_2cf31306[2]),
    .o(al_a7d56e64[10]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_e3d0a508 (
    .a(al_275437c2),
    .b(al_2cf31306[3]),
    .o(al_a7d56e64[11]));
  AL_MAP_LUT5 #(
    .EQN("~(E@D@C@B@A)"),
    .INIT(32'h69969669))
    al_a31c575c (
    .a(al_5411d218),
    .b(al_a7b91d29),
    .c(al_f4b18dcd),
    .d(al_8a6ca59e[6]),
    .e(al_2cf31306[25]),
    .o(al_4c9c0764));
  AL_MAP_LUT3 #(
    .EQN("(C@(B*~A))"),
    .INIT(8'hb4))
    al_5c94036c (
    .a(al_4c9c0764),
    .b(al_2a71f823),
    .c(al_2cf31306[4]),
    .o(al_a7d56e64[12]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_b143ccea (
    .a(al_8a6ca59e[5]),
    .b(al_2cf31306[26]),
    .o(al_f4b18dcd));
  AL_MAP_LUT4 #(
    .EQN("(D@C@B@A)"),
    .INIT(16'h6996))
    al_6dfdfb86 (
    .a(al_8a6ca59e[1]),
    .b(al_8a6ca59e[2]),
    .c(al_2cf31306[29]),
    .d(al_2cf31306[30]),
    .o(al_bfb14c0f));
  AL_MAP_LUT6 #(
    .EQN("(F@(E*(D@C@B@A)))"),
    .INIT(64'h9669ffff69960000))
    al_c4a071e5 (
    .a(al_219561f),
    .b(al_bfb14c0f),
    .c(al_e30f13e9),
    .d(al_f4b18dcd),
    .e(al_2a71f823),
    .f(al_2cf31306[5]),
    .o(al_a7d56e64[13]));
  AL_MAP_LUT3 #(
    .EQN("(C@B@A)"),
    .INIT(8'h96))
    al_e99ad987 (
    .a(al_e30f13e9),
    .b(al_8a6ca59e[3]),
    .c(al_2cf31306[28]),
    .o(al_54bdd1be));
  AL_MAP_LUT5 #(
    .EQN("(E@(D*~(C@B@A)))"),
    .INIT(32'h96ff6900))
    al_720d5e53 (
    .a(al_b130642e[0]),
    .b(al_54bdd1be),
    .c(al_f4b18dcd),
    .d(al_2a71f823),
    .e(al_2cf31306[6]),
    .o(al_a7d56e64[14]));
  AL_MAP_LUT5 #(
    .EQN("(E@(D*(C@B@A)))"),
    .INIT(32'h69ff9600))
    al_fe465bf0 (
    .a(al_a7b91d29),
    .b(al_e30f13e9),
    .c(al_3d188dba),
    .d(al_2a71f823),
    .e(al_2cf31306[7]),
    .o(al_a7d56e64[15]));
  AL_MAP_LUT5 #(
    .EQN("(D@(B*~(E@C@A)))"),
    .INIT(32'hb7487b84))
    al_638ca3f3 (
    .a(al_a7b91d29),
    .b(al_2a71f823),
    .c(al_8a6ca59e[7]),
    .d(al_2cf31306[8]),
    .e(al_2cf31306[24]),
    .o(al_a7d56e64[16]));
  AL_MAP_LUT5 #(
    .EQN("(D@(B*~(E@C@A)))"),
    .INIT(32'hb7487b84))
    al_b3736838 (
    .a(al_bfb14c0f),
    .b(al_2a71f823),
    .c(al_8a6ca59e[6]),
    .d(al_2cf31306[9]),
    .e(al_2cf31306[25]),
    .o(al_a7d56e64[17]));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*~(B@A)))"),
    .INIT(16'h6f90))
    al_f6de39ad (
    .a(al_b130642e[0]),
    .b(al_f4b18dcd),
    .c(al_2a71f823),
    .d(al_2cf31306[10]),
    .o(al_a7d56e64[18]));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*(B@A)))"),
    .INIT(16'h9f60))
    al_8853877b (
    .a(al_e30f13e9),
    .b(al_3d188dba),
    .c(al_2a71f823),
    .d(al_2cf31306[11]),
    .o(al_a7d56e64[19]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_d59bf2 (
    .a(al_4fb560ef),
    .b(al_2a71f823),
    .c(al_8a6ca59e[1]),
    .o(al_a7d56e64[1]));
  AL_MAP_LUT4 #(
    .EQN("(C@(A*~(D@B)))"),
    .INIT(16'h78d2))
    al_c4258b4 (
    .a(al_2a71f823),
    .b(al_8a6ca59e[3]),
    .c(al_2cf31306[12]),
    .d(al_2cf31306[28]),
    .o(al_a7d56e64[20]));
  AL_MAP_LUT4 #(
    .EQN("(C@(A*~(D@B)))"),
    .INIT(16'h78d2))
    al_ceeee258 (
    .a(al_2a71f823),
    .b(al_8a6ca59e[2]),
    .c(al_2cf31306[13]),
    .d(al_2cf31306[29]),
    .o(al_a7d56e64[21]));
  AL_MAP_LUT4 #(
    .EQN("(C@(A*~(D@B)))"),
    .INIT(16'h78d2))
    al_461b38bd (
    .a(al_2a71f823),
    .b(al_8a6ca59e[7]),
    .c(al_2cf31306[14]),
    .d(al_2cf31306[24]),
    .o(al_a7d56e64[22]));
  AL_MAP_LUT5 #(
    .EQN("(D@(B*~(E@C@A)))"),
    .INIT(32'hb7487b84))
    al_c9d6ce01 (
    .a(al_5411d218),
    .b(al_2a71f823),
    .c(al_8a6ca59e[6]),
    .d(al_2cf31306[15]),
    .e(al_2cf31306[25]),
    .o(al_a7d56e64[23]));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*~(B@A)))"),
    .INIT(16'h6f90))
    al_9b2667b (
    .a(al_219561f),
    .b(al_f4b18dcd),
    .c(al_2a71f823),
    .d(al_2cf31306[16]),
    .o(al_a7d56e64[24]));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*(B@A)))"),
    .INIT(16'h9f60))
    al_1924ecd4 (
    .a(al_e30f13e9),
    .b(al_f4b18dcd),
    .c(al_2a71f823),
    .d(al_2cf31306[17]),
    .o(al_a7d56e64[25]));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*(B@A)))"),
    .INIT(16'h9f60))
    al_11baff80 (
    .a(al_54bdd1be),
    .b(al_5411d218),
    .c(al_2a71f823),
    .d(al_2cf31306[18]),
    .o(al_a7d56e64[26]));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*(B@A)))"),
    .INIT(16'h9f60))
    al_62b400f6 (
    .a(al_219561f),
    .b(al_a7b91d29),
    .c(al_2a71f823),
    .d(al_2cf31306[19]),
    .o(al_a7d56e64[27]));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*~(B@A)))"),
    .INIT(16'h6f90))
    al_a88f48bf (
    .a(al_bfb14c0f),
    .b(al_f4b18dcd),
    .c(al_2a71f823),
    .d(al_2cf31306[20]),
    .o(al_a7d56e64[28]));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*~(B@A)))"),
    .INIT(16'h6f90))
    al_2ffb6df8 (
    .a(al_b130642e[0]),
    .b(al_e30f13e9),
    .c(al_2a71f823),
    .d(al_2cf31306[21]),
    .o(al_a7d56e64[29]));
  AL_MAP_LUT4 #(
    .EQN("(D*~((B@A))*~(C)+D*(B@A)*~(C)+~(D)*(B@A)*C+D*(B@A)*C)"),
    .INIT(16'h6f60))
    al_5a378330 (
    .a(al_4fb560ef),
    .b(al_f4b18dcd),
    .c(al_2a71f823),
    .d(al_8a6ca59e[2]),
    .o(al_a7d56e64[2]));
  AL_MAP_LUT5 #(
    .EQN("(D@(B*(E@C@A)))"),
    .INIT(32'h7b84b748))
    al_af5e5c8b (
    .a(al_3d188dba),
    .b(al_2a71f823),
    .c(al_8a6ca59e[3]),
    .d(al_2cf31306[22]),
    .e(al_2cf31306[28]),
    .o(al_a7d56e64[30]));
  AL_MAP_LUT4 #(
    .EQN("(C@(A*~(D@B)))"),
    .INIT(16'h78d2))
    al_bb9c8e9c (
    .a(al_2a71f823),
    .b(al_8a6ca59e[2]),
    .c(al_2cf31306[23]),
    .d(al_2cf31306[29]),
    .o(al_a7d56e64[31]));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~((C@B@A))*~(D)+~E*(C@B@A)*~(D)+~(~E)*(C@B@A)*D+~E*(C@B@A)*D)"),
    .INIT(32'h69ff6900))
    al_34ea70dd (
    .a(al_219561f),
    .b(al_e30f13e9),
    .c(al_f4b18dcd),
    .d(al_2a71f823),
    .e(al_8a6ca59e[3]),
    .o(al_a7d56e64[3]));
  AL_MAP_LUT5 #(
    .EQN("(E*~((C@B@A))*~(D)+E*(C@B@A)*~(D)+~(E)*(C@B@A)*D+E*(C@B@A)*D)"),
    .INIT(32'h96ff9600))
    al_c7e8f8f6 (
    .a(al_54bdd1be),
    .b(al_5411d218),
    .c(al_f4b18dcd),
    .d(al_2a71f823),
    .e(al_8a6ca59e[4]),
    .o(al_a7d56e64[4]));
  AL_MAP_LUT4 #(
    .EQN("(D@C@B@A)"),
    .INIT(16'h6996))
    al_87ed432f (
    .a(al_8a6ca59e[1]),
    .b(al_8a6ca59e[7]),
    .c(al_2cf31306[24]),
    .d(al_2cf31306[30]),
    .o(al_5411d218));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_63b65d75 (
    .a(al_219561f),
    .b(al_5411d218),
    .o(al_4fb560ef));
  AL_MAP_LUT5 #(
    .EQN("(E*~((C@B@A))*~(D)+E*(C@B@A)*~(D)+~(E)*(C@B@A)*D+E*(C@B@A)*D)"),
    .INIT(32'h96ff9600))
    al_57989698 (
    .a(al_4fb560ef),
    .b(al_a7b91d29),
    .c(al_e30f13e9),
    .d(al_2a71f823),
    .e(al_8a6ca59e[5]),
    .o(al_a7d56e64[5]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_4a195ea9 (
    .a(al_8a6ca59e[4]),
    .b(al_2cf31306[27]),
    .o(al_e30f13e9));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_d62ea490 (
    .a(al_8a6ca59e[0]),
    .b(al_2cf31306[31]),
    .o(al_3d188dba));
  AL_MAP_LUT4 #(
    .EQN("(D@C@B@A)"),
    .INIT(16'h6996))
    al_a941f1b3 (
    .a(al_8a6ca59e[2]),
    .b(al_8a6ca59e[3]),
    .c(al_2cf31306[28]),
    .d(al_2cf31306[29]),
    .o(al_a7b91d29));
  AL_MAP_LUT3 #(
    .EQN("(C@B@A)"),
    .INIT(8'h96))
    al_cbe2681e (
    .a(al_3d188dba),
    .b(al_8a6ca59e[6]),
    .c(al_2cf31306[25]),
    .o(al_219561f));
  AL_MAP_LUT3 #(
    .EQN("(C@B@A)"),
    .INIT(8'h96))
    al_c590e72d (
    .a(al_3d188dba),
    .b(al_8a6ca59e[1]),
    .c(al_2cf31306[30]),
    .o(al_b130642e[0]));
  AL_MAP_LUT6 #(
    .EQN("(E@(D*~(F@C@B@A)))"),
    .INIT(64'h69ff960096ff6900))
    al_25f8ae63 (
    .a(al_b130642e[0]),
    .b(al_a7b91d29),
    .c(al_f4b18dcd),
    .d(al_2a71f823),
    .e(al_8a6ca59e[6]),
    .f(al_2cf31306[25]),
    .o(al_a7d56e64[6]));
  AL_MAP_LUT6 #(
    .EQN("~(F@E@D@C@B@A)"),
    .INIT(64'h9669699669969669))
    al_25919cc7 (
    .a(al_e30f13e9),
    .b(al_f4b18dcd),
    .c(al_8a6ca59e[2]),
    .d(al_8a6ca59e[7]),
    .e(al_2cf31306[24]),
    .f(al_2cf31306[29]),
    .o(al_c78fe3c1));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~((B@A))*~(C)+~D*(B@A)*~(C)+~(~D)*(B@A)*C+~D*(B@A)*C)"),
    .INIT(16'h9f90))
    al_524fadcf (
    .a(al_c78fe3c1),
    .b(al_3d188dba),
    .c(al_2a71f823),
    .d(al_8a6ca59e[7]),
    .o(al_a7d56e64[7]));
  AL_MAP_LUT6 #(
    .EQN("(B*(F@E@D@C@A))"),
    .INIT(64'h8448488448848448))
    al_91a04c6b (
    .a(al_54bdd1be),
    .b(al_2a71f823),
    .c(al_8a6ca59e[6]),
    .d(al_8a6ca59e[7]),
    .e(al_2cf31306[24]),
    .f(al_2cf31306[25]),
    .o(al_275437c2));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_9502c298 (
    .a(al_275437c2),
    .b(al_2cf31306[0]),
    .o(al_a7d56e64[8]));
  AL_MAP_LUT6 #(
    .EQN("(E@(C*(F@D@B@A)))"),
    .INIT(64'h9f6f60906f9f9060))
    al_7c3957ee (
    .a(al_a7b91d29),
    .b(al_f4b18dcd),
    .c(al_2a71f823),
    .d(al_8a6ca59e[6]),
    .e(al_2cf31306[1]),
    .f(al_2cf31306[25]),
    .o(al_a7d56e64[9]));
  AL_DFF_X al_8e787e71 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a7d56e64[0]),
    .en(tx_clk_en),
    .sr(al_48fcd383[2]),
    .ss(1'b0),
    .q(al_2cf31306[0]));
  AL_DFF_X al_ee7fdb39 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a7d56e64[9]),
    .en(tx_clk_en),
    .sr(al_48fcd383[2]),
    .ss(1'b0),
    .q(al_2cf31306[9]));
  AL_DFF_X al_3e8c5e65 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a7d56e64[10]),
    .en(tx_clk_en),
    .sr(al_48fcd383[2]),
    .ss(1'b0),
    .q(al_2cf31306[10]));
  AL_DFF_X al_3e477b36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a7d56e64[11]),
    .en(tx_clk_en),
    .sr(al_48fcd383[2]),
    .ss(1'b0),
    .q(al_2cf31306[11]));
  AL_DFF_X al_858a0e95 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a7d56e64[12]),
    .en(tx_clk_en),
    .sr(al_48fcd383[2]),
    .ss(1'b0),
    .q(al_2cf31306[12]));
  AL_DFF_X al_d3b0a930 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a7d56e64[13]),
    .en(tx_clk_en),
    .sr(al_48fcd383[2]),
    .ss(1'b0),
    .q(al_2cf31306[13]));
  AL_DFF_X al_e4e63ab7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a7d56e64[14]),
    .en(tx_clk_en),
    .sr(al_48fcd383[2]),
    .ss(1'b0),
    .q(al_2cf31306[14]));
  AL_DFF_X al_b09582d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a7d56e64[15]),
    .en(tx_clk_en),
    .sr(al_48fcd383[2]),
    .ss(1'b0),
    .q(al_2cf31306[15]));
  AL_DFF_X al_5150b17f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a7d56e64[16]),
    .en(tx_clk_en),
    .sr(al_48fcd383[2]),
    .ss(1'b0),
    .q(al_2cf31306[16]));
  AL_DFF_X al_73a764e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a7d56e64[17]),
    .en(tx_clk_en),
    .sr(al_48fcd383[2]),
    .ss(1'b0),
    .q(al_2cf31306[17]));
  AL_DFF_X al_1eb83e66 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a7d56e64[18]),
    .en(tx_clk_en),
    .sr(al_48fcd383[2]),
    .ss(1'b0),
    .q(al_2cf31306[18]));
  AL_DFF_X al_d397d3b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a7d56e64[1]),
    .en(tx_clk_en),
    .sr(al_48fcd383[2]),
    .ss(1'b0),
    .q(al_2cf31306[1]));
  AL_DFF_X al_792c6fb7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a7d56e64[19]),
    .en(tx_clk_en),
    .sr(al_48fcd383[2]),
    .ss(1'b0),
    .q(al_2cf31306[19]));
  AL_DFF_X al_e1da6a12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a7d56e64[20]),
    .en(tx_clk_en),
    .sr(al_48fcd383[2]),
    .ss(1'b0),
    .q(al_2cf31306[20]));
  AL_DFF_X al_9d5c2a3d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a7d56e64[21]),
    .en(tx_clk_en),
    .sr(al_48fcd383[2]),
    .ss(1'b0),
    .q(al_2cf31306[21]));
  AL_DFF_X al_96af2aca (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a7d56e64[22]),
    .en(tx_clk_en),
    .sr(al_48fcd383[2]),
    .ss(1'b0),
    .q(al_2cf31306[22]));
  AL_DFF_X al_90cfeab9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a7d56e64[23]),
    .en(tx_clk_en),
    .sr(al_48fcd383[2]),
    .ss(1'b0),
    .q(al_2cf31306[23]));
  AL_DFF_X al_505a5c4f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a7d56e64[24]),
    .en(tx_clk_en),
    .sr(al_48fcd383[2]),
    .ss(1'b0),
    .q(al_2cf31306[24]));
  AL_DFF_X al_24194b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a7d56e64[25]),
    .en(tx_clk_en),
    .sr(al_48fcd383[2]),
    .ss(1'b0),
    .q(al_2cf31306[25]));
  AL_DFF_X al_7d1f3a58 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a7d56e64[26]),
    .en(tx_clk_en),
    .sr(al_48fcd383[2]),
    .ss(1'b0),
    .q(al_2cf31306[26]));
  AL_DFF_X al_5ba87b62 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a7d56e64[27]),
    .en(tx_clk_en),
    .sr(al_48fcd383[2]),
    .ss(1'b0),
    .q(al_2cf31306[27]));
  AL_DFF_X al_6c5c23e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a7d56e64[28]),
    .en(tx_clk_en),
    .sr(al_48fcd383[2]),
    .ss(1'b0),
    .q(al_2cf31306[28]));
  AL_DFF_X al_8d531918 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a7d56e64[2]),
    .en(tx_clk_en),
    .sr(al_48fcd383[2]),
    .ss(1'b0),
    .q(al_2cf31306[2]));
  AL_DFF_X al_1b62185d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a7d56e64[29]),
    .en(tx_clk_en),
    .sr(al_48fcd383[2]),
    .ss(1'b0),
    .q(al_2cf31306[29]));
  AL_DFF_X al_b120568a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a7d56e64[30]),
    .en(tx_clk_en),
    .sr(al_48fcd383[2]),
    .ss(1'b0),
    .q(al_2cf31306[30]));
  AL_DFF_X al_baa32a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a7d56e64[31]),
    .en(tx_clk_en),
    .sr(al_48fcd383[2]),
    .ss(1'b0),
    .q(al_2cf31306[31]));
  AL_DFF_X al_e17f306c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a7d56e64[3]),
    .en(tx_clk_en),
    .sr(al_48fcd383[2]),
    .ss(1'b0),
    .q(al_2cf31306[3]));
  AL_DFF_X al_f38c789a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a7d56e64[4]),
    .en(tx_clk_en),
    .sr(al_48fcd383[2]),
    .ss(1'b0),
    .q(al_2cf31306[4]));
  AL_DFF_X al_3233e361 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a7d56e64[5]),
    .en(tx_clk_en),
    .sr(al_48fcd383[2]),
    .ss(1'b0),
    .q(al_2cf31306[5]));
  AL_DFF_X al_d169b1ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a7d56e64[6]),
    .en(tx_clk_en),
    .sr(al_48fcd383[2]),
    .ss(1'b0),
    .q(al_2cf31306[6]));
  AL_DFF_X al_ecabd58a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a7d56e64[7]),
    .en(tx_clk_en),
    .sr(al_48fcd383[2]),
    .ss(1'b0),
    .q(al_2cf31306[7]));
  AL_DFF_X al_31274d4f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a7d56e64[8]),
    .en(tx_clk_en),
    .sr(al_48fcd383[2]),
    .ss(1'b0),
    .q(al_2cf31306[8]));
  AL_DFF_X al_7d62b7cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b3c5207a),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_2a71f823));
  AL_DFF_X al_3ba766bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_964d579),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_e396ca5d));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_7cbd1c9d (
    .a(al_cbafc250),
    .b(al_8a6ca59e[0]),
    .o(al_f83013e9[0]));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~A)*~(D)*~(B)+~(~C*~A)*D*~(B)+~(~(~C*~A))*D*B+~(~C*~A)*D*B)"),
    .INIT(16'hfe32))
    al_b5b07600 (
    .a(al_f83013e9[0]),
    .b(al_e396ca5d),
    .c(al_d75651de),
    .d(al_2cf31306[31]),
    .o(al_96e5a141[0]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_7c3e9c1 (
    .a(al_cbafc250),
    .b(al_8a6ca59e[1]),
    .o(al_f83013e9[1]));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~A)*~(D)*~(B)+~(~C*~A)*D*~(B)+~(~(~C*~A))*D*B+~(~C*~A)*D*B)"),
    .INIT(16'hfe32))
    al_f97b7429 (
    .a(al_f83013e9[1]),
    .b(al_e396ca5d),
    .c(al_d75651de),
    .d(al_2cf31306[30]),
    .o(al_96e5a141[1]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_94c64f9d (
    .a(al_cbafc250),
    .b(al_8a6ca59e[2]),
    .o(al_f83013e9[2]));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~A)*~(D)*~(B)+~(~C*~A)*D*~(B)+~(~(~C*~A))*D*B+~(~C*~A)*D*B)"),
    .INIT(16'hfe32))
    al_178c641d (
    .a(al_f83013e9[2]),
    .b(al_e396ca5d),
    .c(al_d75651de),
    .d(al_2cf31306[29]),
    .o(al_96e5a141[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_dd658972 (
    .a(al_cbafc250),
    .b(al_8a6ca59e[3]),
    .o(al_f83013e9[3]));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~A)*~(D)*~(B)+~(~C*~A)*D*~(B)+~(~(~C*~A))*D*B+~(~C*~A)*D*B)"),
    .INIT(16'hfe32))
    al_ea11ad56 (
    .a(al_f83013e9[3]),
    .b(al_e396ca5d),
    .c(al_d75651de),
    .d(al_2cf31306[28]),
    .o(al_96e5a141[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_b87e4624 (
    .a(al_cbafc250),
    .b(al_8a6ca59e[4]),
    .o(al_f83013e9[4]));
  AL_MAP_LUT4 #(
    .EQN("((~C*A)*~(D)*~(B)+(~C*A)*D*~(B)+~((~C*A))*D*B+(~C*A)*D*B)"),
    .INIT(16'hce02))
    al_51c8968e (
    .a(al_f83013e9[4]),
    .b(al_e396ca5d),
    .c(al_d75651de),
    .d(al_2cf31306[27]),
    .o(al_96e5a141[4]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_8b9c90c5 (
    .a(al_cbafc250),
    .b(al_8a6ca59e[5]),
    .o(al_f83013e9[5]));
  AL_MAP_LUT4 #(
    .EQN("((~C*A)*~(D)*~(B)+(~C*A)*D*~(B)+~((~C*A))*D*B+(~C*A)*D*B)"),
    .INIT(16'hce02))
    al_52d061ff (
    .a(al_f83013e9[5]),
    .b(al_e396ca5d),
    .c(al_d75651de),
    .d(al_2cf31306[26]),
    .o(al_96e5a141[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_b05675d5 (
    .a(al_cbafc250),
    .b(al_8a6ca59e[6]),
    .o(al_f83013e9[6]));
  AL_MAP_LUT4 #(
    .EQN("((~C*A)*~(D)*~(B)+(~C*A)*D*~(B)+~((~C*A))*D*B+(~C*A)*D*B)"),
    .INIT(16'hce02))
    al_fa558d1e (
    .a(al_f83013e9[6]),
    .b(al_e396ca5d),
    .c(al_d75651de),
    .d(al_2cf31306[25]),
    .o(al_96e5a141[6]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_6ef9c77e (
    .a(al_cbafc250),
    .b(al_8a6ca59e[7]),
    .o(al_f83013e9[7]));
  AL_MAP_LUT4 #(
    .EQN("((~C*A)*~(D)*~(B)+(~C*A)*D*~(B)+~((~C*A))*D*B+(~C*A)*D*B)"),
    .INIT(16'hce02))
    al_6111f5a1 (
    .a(al_f83013e9[7]),
    .b(al_e396ca5d),
    .c(al_d75651de),
    .d(al_2cf31306[24]),
    .o(al_96e5a141[7]));
  AL_DFF_X al_5737c9dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1491ad5),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_7cd73f8f));
  AL_DFF_X al_8c4924c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5c023966),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1bfb1d64));
  AL_MAP_LUT6 #(
    .EQN("(~C*(F*~((E*D*A))*~(B)+F*(E*D*A)*~(B)+~(F)*(E*D*A)*B+F*(E*D*A)*B))"),
    .INIT(64'h0b03030308000000))
    al_4fe0d5 (
    .a(al_2179357c),
    .b(al_5d1a6fb0),
    .c(al_6b4499fc),
    .d(al_64e175a6),
    .e(al_e00c8785[0]),
    .f(al_1bfb1d64),
    .o(al_5c023966));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_d826c9da (
    .a(tx_clk_en),
    .b(al_48fcd383[4]),
    .o(al_5d1a6fb0));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_a30e4a33 (
    .a(al_e00c8785[1]),
    .b(al_e00c8785[2]),
    .c(al_e00c8785[3]),
    .d(al_e00c8785[4]),
    .o(al_44998c84));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_ab71f10b (
    .a(al_44998c84),
    .b(al_e00c8785[5]),
    .c(al_e00c8785[6]),
    .d(al_e00c8785[7]),
    .o(al_2179357c));
  AL_DFF_X al_6ae0c7c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_76966ac9),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_af1ac2b6));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*A)"),
    .INIT(64'h8000000000000000))
    al_5c42d058 (
    .a(al_8a6ca59e[2]),
    .b(al_8a6ca59e[3]),
    .c(al_8a6ca59e[4]),
    .d(al_8a6ca59e[5]),
    .e(al_8a6ca59e[6]),
    .f(al_8a6ca59e[7]),
    .o(al_4f8a4577));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_e9a0d5f2 (
    .a(al_4f8a4577),
    .b(al_64e175a6),
    .c(al_8a6ca59e[0]),
    .d(al_8a6ca59e[1]),
    .o(al_bca5d36c));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT(16'h0b08))
    al_a0141f7 (
    .a(al_bca5d36c),
    .b(al_5d1a6fb0),
    .c(al_6b4499fc),
    .d(al_af1ac2b6),
    .o(al_76966ac9));
  AL_DFF_X al_a42b90cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ca9e38f4),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_75182ad3));
  AL_MAP_LUT6 #(
    .EQN("(~C*(F*~((E*D*A))*~(B)+F*(E*D*A)*~(B)+~(F)*(E*D*A)*B+F*(E*D*A)*B))"),
    .INIT(64'h0b03030308000000))
    al_3a94dac2 (
    .a(al_bbe3a962),
    .b(al_5d1a6fb0),
    .c(al_6b4499fc),
    .d(al_64e175a6),
    .e(al_84c0beb4[0]),
    .f(al_75182ad3),
    .o(al_ca9e38f4));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_e88d9668 (
    .a(al_84c0beb4[1]),
    .b(al_84c0beb4[2]),
    .c(al_84c0beb4[3]),
    .d(al_84c0beb4[4]),
    .o(al_f7494ece));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_1d8692e4 (
    .a(al_f7494ece),
    .b(al_84c0beb4[5]),
    .c(al_84c0beb4[6]),
    .d(al_84c0beb4[7]),
    .o(al_bbe3a962));
  AL_DFF_X al_ad8bcc05 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_54fc2cdd),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5ad7d7e7));
  AL_MAP_LUT6 #(
    .EQN("(~C*(F*~((E*D*A))*~(B)+F*(E*D*A)*~(B)+~(F)*(E*D*A)*B+F*(E*D*A)*B))"),
    .INIT(64'h0b03030308000000))
    al_b96b7292 (
    .a(al_65b028e9),
    .b(al_5d1a6fb0),
    .c(al_6b4499fc),
    .d(al_64e175a6),
    .e(al_9affd881[0]),
    .f(al_5ad7d7e7),
    .o(al_54fc2cdd));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_5a327671 (
    .a(al_9affd881[1]),
    .b(al_9affd881[2]),
    .c(al_9affd881[3]),
    .d(al_9affd881[4]),
    .o(al_6300b493));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_9a0c8fb1 (
    .a(al_6300b493),
    .b(al_9affd881[5]),
    .c(al_9affd881[6]),
    .d(al_9affd881[7]),
    .o(al_65b028e9));
  AL_DFF_X al_2dda4e26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c981d7f0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c5664b3b));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*A)"),
    .INIT(64'h8000000000000000))
    al_5799c7b4 (
    .a(al_64e175a6),
    .b(al_4d46dbf7[0]),
    .c(al_4d46dbf7[1]),
    .d(al_4d46dbf7[2]),
    .e(al_4d46dbf7[3]),
    .f(al_4d46dbf7[4]),
    .o(al_1ce38576));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_db5a6450 (
    .a(al_1ce38576),
    .b(al_4d46dbf7[5]),
    .c(al_4d46dbf7[6]),
    .d(al_4d46dbf7[7]),
    .o(al_7c03a443));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT(16'h0b08))
    al_1dc4e0b (
    .a(al_7c03a443),
    .b(al_5d1a6fb0),
    .c(al_6b4499fc),
    .d(al_c5664b3b),
    .o(al_c981d7f0));
  AL_DFF_X al_ac0bd0d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d5243429),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9f6ea2ef));
  AL_MAP_LUT5 #(
    .EQN("(~C*(E*~(A)*~((D*B))+E*A*~((D*B))+~(E)*A*(D*B)+E*A*(D*B)))"),
    .INIT(32'h0b0f0800))
    al_adc76e28 (
    .a(al_7c03a443),
    .b(tx_clk_en),
    .c(al_6b4499fc),
    .d(al_48fcd383[5]),
    .e(al_9f6ea2ef),
    .o(al_d5243429));
  AL_DFF_X al_2d42802e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5f85f29c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad4aba0));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h3120))
    al_2b3294c9 (
    .a(al_5d1a6fb0),
    .b(al_6b4499fc),
    .c(al_e00c8785[0]),
    .d(al_ad4aba0),
    .o(al_5f85f29c));
  AL_DFF_X al_3eecc52 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cf06a90),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_c52cf3e8));
  AL_DFF_X al_d7421c6b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4421c6bd),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_6fa8f988));
  AL_DFF_X al_d9775949 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4be4ecdd),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_20a6f635));
  AL_DFF_X al_5cd8ec3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f192c825),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_5b769262));
  AL_DFF_X al_989f6200 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_17387d1),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_548d2e8d));
  AL_DFF_X al_c220aa3f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9f207ad1),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_ee3bb963));
  AL_DFF_X al_908722eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4973ef09),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_1f6fed00));
  AL_DFF_X al_9cb992bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_85bba154),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_b7729dd8));
  AL_DFF_X al_cd281a4c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1d84107f),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_85bba154));
  AL_DFF_X al_c361ba4b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_114ce5a4),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_c35ead5c));
  AL_DFF_X al_f60d5c07 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c59c6deb),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_ea30f787));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_6ed832a1 (
    .a(al_183e87f4[0]),
    .b(al_64fd2ef5[0]),
    .c(al_af6614da),
    .o(al_24da7d44[0]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_27ed91a9 (
    .a(al_183e87f4[10]),
    .b(al_64fd2ef5[10]),
    .c(al_af6614da),
    .o(al_24da7d44[10]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_7a180426 (
    .a(al_183e87f4[11]),
    .b(al_64fd2ef5[11]),
    .c(al_af6614da),
    .o(al_24da7d44[11]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_25d0c11f (
    .a(al_183e87f4[12]),
    .b(al_64fd2ef5[12]),
    .c(al_af6614da),
    .o(al_24da7d44[12]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_c53abdf2 (
    .a(al_183e87f4[13]),
    .b(al_64fd2ef5[13]),
    .c(al_af6614da),
    .o(al_24da7d44[13]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_19f6345b (
    .a(al_183e87f4[1]),
    .b(al_64fd2ef5[1]),
    .c(al_af6614da),
    .o(al_24da7d44[1]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_752258a0 (
    .a(al_183e87f4[2]),
    .b(al_64fd2ef5[2]),
    .c(al_af6614da),
    .o(al_24da7d44[2]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_69d2743d (
    .a(al_183e87f4[3]),
    .b(al_64fd2ef5[3]),
    .c(al_af6614da),
    .o(al_24da7d44[3]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_c9489a6b (
    .a(al_183e87f4[4]),
    .b(al_64fd2ef5[4]),
    .c(al_af6614da),
    .o(al_24da7d44[4]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_8c9beb18 (
    .a(al_183e87f4[5]),
    .b(al_64fd2ef5[5]),
    .c(al_af6614da),
    .o(al_24da7d44[5]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_c7827c6f (
    .a(al_183e87f4[6]),
    .b(al_64fd2ef5[6]),
    .c(al_af6614da),
    .o(al_24da7d44[6]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_531797ab (
    .a(al_183e87f4[7]),
    .b(al_64fd2ef5[7]),
    .c(al_af6614da),
    .o(al_24da7d44[7]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_151c7a9f (
    .a(al_183e87f4[8]),
    .b(al_64fd2ef5[8]),
    .c(al_af6614da),
    .o(al_24da7d44[8]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d977584 (
    .a(al_183e87f4[9]),
    .b(al_64fd2ef5[9]),
    .c(al_af6614da),
    .o(al_24da7d44[9]));
  AL_DFF_X al_787ea2b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_7ac4c27f),
    .en(al_520be21e),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_af6614da));
  AL_DFF_X al_7915f0c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_397de144),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_d75651de));
  AL_DFF_X al_fbd60f69 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ec9f94d8),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1e17be4));
  AL_MAP_LUT6 #(
    .EQN("(~B*(D*~(C)*~((~(~F*~E)*A))+D*C*~((~(~F*~E)*A))+~(D)*C*(~(~F*~E)*A)+D*C*(~(~F*~E)*A)))"),
    .INIT(64'h3120312031203300))
    al_e9e73cd3 (
    .a(tx_clk_en),
    .b(al_6b4499fc),
    .c(al_10fc4c0e),
    .d(al_d1e17be4),
    .e(al_a494216e),
    .f(al_33f2071f),
    .o(al_ec9f94d8));
  AL_DFF_X al_a8d19d62 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_dd9e938b),
    .en(al_520be21e),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_d3482891));
  AL_DFF_X al_a3332f23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_8cc75feb),
    .en(al_520be21e),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_ea441981));
  AL_DFF_X al_1c376cd3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_643ac1f2),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_cf085f09));
  AL_DFF_X al_a2295bf5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a6c89001),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_f6643499));
  AL_DFF_X al_30417ce8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_54081406),
    .en(al_520be21e),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_edc29fee));
  AL_DFF_X al_9d18d43d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_a1a0ec14),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_206f470e));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    al_22b57374 (
    .a(al_a140f198),
    .b(al_bff87853[0]),
    .c(al_bff87853[3]),
    .d(al_bff87853[11]),
    .o(al_f92f3a06));
  AL_DFF_X al_23581d37 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_47e79db6),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e175a6));
  AL_MAP_LUT6 #(
    .EQN("(~C*(E*~((~F*A))*~((D*B))+E*(~F*A)*~((D*B))+~(E)*(~F*A)*(D*B)+E*(~F*A)*(D*B)))"),
    .INIT(64'h030f00000b0f0800))
    al_7d12c227 (
    .a(al_2337d80f),
    .b(tx_clk_en),
    .c(al_6b4499fc),
    .d(al_177c7491),
    .e(al_64e175a6),
    .f(al_21d722fe),
    .o(al_47e79db6));
  AL_DFF_X al_1890dfe9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e03ae0c1),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_3475fb1c));
  AL_DFF_X al_4d9486ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_508b6c4c),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_8b86ece7));
  AL_DFF_X al_1a5e3d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_66382828),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_4dac203f));
  AL_DFF_X al_d20954e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5156ba29),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_6980bc30));
  AL_DFF_X al_99b1a37e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_8aeddbc),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_2b1074ba));
  AL_DFF_X al_a97c3acf (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_95d27a4c),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_b65fd623));
  AL_DFF_X al_fe145f59 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ab82ee9a),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_21d722fe));
  AL_DFF_X al_c58ed4da (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_6b5283b3),
    .en(al_520be21e),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_f731da11));
  AL_DFF_X al_cc635404 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_8f030415),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_cbafc250));
  AL_DFF_X al_a3c47b1e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_6b2f12fa),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_3e886516));
  AL_DFF_X al_5afb9a6a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_bb3ef93c),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_e199650d));
  AL_DFF_X al_743699e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ffd3f5d1),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_643ac1f2));
  AL_DFF_X al_cf1af11a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_da8b063f),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_fdd1f60e));
  AL_DFF_X al_e316e1db (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_70a59d2e),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_642e830e));
  AL_DFF_X al_6cfd9ec2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f2d6f40b),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_4a548f7c));
  AL_DFF_X al_8efdc5fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e5fcf9b1),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_f2f960a1));
  AL_DFF_X al_5288e35b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4e7d0870),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_e5fcf9b1));
  AL_DFF_X al_12b68c12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_db73eae9),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_eb5c4882));
  AL_DFF_X al_a2c9ce3a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_64c768d),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_33f2071f));
  AL_DFF_X al_ce0917ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4854aa2f),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_a978a29f));
  AL_DFF_X al_cf825408 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(gmii_col),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_d27166fa));
  AL_DFF_X al_930bc316 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_977227b4),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_f92026f1));
  AL_DFF_X al_d9776907 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2337d80f),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9a8c459a));
  AL_DFF_X al_8e9f7b45 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4d4a65fe),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_d224660a));
  AL_DFF_X al_700c8006 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_7ffb8465),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_6490a8fc));
  AL_DFF_X al_8fea456d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e1420a1f),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_f52ae365));
  AL_DFF_X al_9ba52cac (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_eb5c4882),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_b348c1a2));
  AL_DFF_X al_93d93e76 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_72403be8),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_be1d3817));
  AL_DFF_X al_2f05a0a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_7f7f4148),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_f28e4921));
  AL_DFF_X al_36f0c899 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f92f3a06),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_4b2213d6));
  AL_DFF_X al_429ade15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_1a7bad30),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_3620963e));
  AL_DFF_X al_6d02c1d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e5091a32),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_b1328a1f));
  AL_DFF_X al_ea4464c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_98e25f8d),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_72403be8));
  AL_DFF_X al_42596519 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4a89f542),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_bea385e7));
  AL_DFF_X al_7d033d82 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_567fa47e),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(tx_status_vld));
  AL_DFF_X al_8c88e2ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_8b965f41),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_25d4a5f3));
  AL_DFF_X al_7eeb2607 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_aa6ddd9b),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_e2a3cd9));
  AL_DFF_X al_f151ce08 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b0eb70b2),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_c388f857));
  AL_DFF_X al_30e33239 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_56978088),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_6a534a0a));
  AL_DFF_X al_da5ee933 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_6a534a0a),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_4d3e0511));
  AL_DFF_X al_7d08bc32 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e336c621),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_56978088));
  AL_DFF_X al_b1a3f44b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4d7216c9),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_13f48428));
  AL_DFF_X al_a630f64b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_acdc1781),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_177c7491));
  AL_DFF_X al_12b91b95 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_81aa4d04),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_77192586));
  AL_DFF_X al_62b7fded (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_81cdbd25),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_1d8c2b07));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_c7315609 (
    .a(1'b0),
    .o({al_4c385591,open_n14}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_7d6c4b9f (
    .a(al_e512aff[0]),
    .b(1'b1),
    .c(al_4c385591),
    .o({al_3fd7c40d,al_f5f472e[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ff56fdbe (
    .a(al_e512aff[1]),
    .b(1'b0),
    .c(al_3fd7c40d),
    .o({al_cf7c6c77,al_f5f472e[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_7372d416 (
    .a(al_e512aff[2]),
    .b(1'b0),
    .c(al_cf7c6c77),
    .o({al_de861c69,al_f5f472e[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_dad88db4 (
    .a(al_e512aff[3]),
    .b(1'b0),
    .c(al_de861c69),
    .o({al_bf96f833,al_f5f472e[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_8ea6203a (
    .a(al_e512aff[4]),
    .b(1'b0),
    .c(al_bf96f833),
    .o({al_191a34b5,al_f5f472e[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_2cffa80a (
    .a(al_e512aff[5]),
    .b(1'b0),
    .c(al_191a34b5),
    .o({al_8aa62a5b,al_f5f472e[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a5842f3c (
    .a(al_e512aff[6]),
    .b(1'b0),
    .c(al_8aa62a5b),
    .o({al_3329776d,al_f5f472e[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ff80a4bd (
    .a(al_e512aff[7]),
    .b(1'b0),
    .c(al_3329776d),
    .o({al_30bba5ae,al_f5f472e[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_aec7557f (
    .a(al_e512aff[8]),
    .b(1'b0),
    .c(al_30bba5ae),
    .o({al_f246f984,al_f5f472e[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_9026e224 (
    .a(al_e512aff[9]),
    .b(1'b0),
    .c(al_f246f984),
    .o({al_b8c67773,al_f5f472e[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_552b98a5 (
    .a(al_e512aff[10]),
    .b(1'b0),
    .c(al_b8c67773),
    .o({al_8319735a,al_f5f472e[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d115d599 (
    .a(al_e512aff[11]),
    .b(1'b0),
    .c(al_8319735a),
    .o({al_639b4ff6,al_f5f472e[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c4fec682 (
    .a(al_e512aff[12]),
    .b(1'b0),
    .c(al_639b4ff6),
    .o({al_717e3e2b,al_f5f472e[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_bea28a1b (
    .a(al_e512aff[13]),
    .b(1'b0),
    .c(al_717e3e2b),
    .o({al_8afbeabf,al_f5f472e[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_cb011e53 (
    .a(al_e512aff[14]),
    .b(1'b0),
    .c(al_8afbeabf),
    .o({open_n15,al_f5f472e[14]}));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_6e323730 (
    .a(tx_clk_en),
    .b(al_33f2071f),
    .o(al_520be21e));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_563d649f (
    .a(tx_clk_en),
    .b(al_48fcd383[13]),
    .o(al_40a7c639));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*B*A)"),
    .INIT(64'h0000000000000008))
    al_225fbe27 (
    .a(al_1698ebe9),
    .b(tx_clk_en),
    .c(al_5b769262),
    .d(al_20a6f635),
    .e(al_cbafc250),
    .f(al_be1d3817),
    .o(al_fbfd813b));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    al_1325ccf (
    .a(al_12358921),
    .b(al_5b769262),
    .c(al_72403be8),
    .d(al_cbafc250),
    .o(al_8640fd7b));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(D*~C*B))"),
    .INIT(16'haeaa))
    al_34f2a068 (
    .a(al_8640fd7b),
    .b(al_177c7491),
    .c(al_7fe117d0),
    .d(al_643ac1f2),
    .o(al_df015ce6));
  AL_MAP_LUT6 #(
    .EQN("(F*~(~D*~C)*~(~B*~(E*A)))"),
    .INIT(64'heee0ccc000000000))
    al_8acdde7 (
    .a(al_7fe117d0),
    .b(al_12358921),
    .c(al_77f0ddfc[0]),
    .d(al_77f0ddfc[1]),
    .e(al_642e830e),
    .f(al_af6614da),
    .o(al_742c008b));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(~C*B)))"),
    .INIT(16'h00ae))
    al_639b6189 (
    .a(al_742c008b),
    .b(al_5b769262),
    .c(al_72403be8),
    .d(al_cbafc250),
    .o(al_f192c825));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*~A)"),
    .INIT(32'h00000004))
    al_8ba2474c (
    .a(al_85bba154),
    .b(al_72403be8),
    .c(al_13f48428),
    .d(al_cbafc250),
    .e(al_56978088),
    .o(al_29b24aa7));
  AL_MAP_LUT6 #(
    .EQN("~(~A*~(~(~D*~(E*C))*~(B)*~(F)+~(~D*~(E*C))*B*~(F)+~(~(~D*~(E*C)))*B*F+~(~D*~(E*C))*B*F))"),
    .INIT(64'heeeeeeeefffaffaa))
    al_85737ed (
    .a(al_29b24aa7),
    .b(al_36605837),
    .c(al_7fe117d0),
    .d(al_12358921),
    .e(al_642e830e),
    .f(al_af6614da),
    .o(al_98e25f8d));
  AL_MAP_LUT6 #(
    .EQN("~((C*B)*~((A*~(E*D)))*~(F)+(C*B)*(A*~(E*D))*~(F)+~((C*B))*(A*~(E*D))*F+(C*B)*(A*~(E*D))*F)"),
    .INIT(64'hff5555553f3f3f3f))
    al_7842c970 (
    .a(al_36605837),
    .b(al_7fe117d0),
    .c(al_642e830e),
    .d(al_643ac1f2),
    .e(al_68ba43d4),
    .f(al_af6614da),
    .o(al_93b20b44));
  AL_MAP_LUT5 #(
    .EQN("~(A*~(~E*~D*C*B))"),
    .INIT(32'h555555d5))
    al_800e123c (
    .a(al_93b20b44),
    .b(al_1698ebe9),
    .c(al_ee3bb963),
    .d(al_20a6f635),
    .e(al_cbafc250),
    .o(al_9f207ad1));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_e9baa5ce (
    .a(al_5b769262),
    .b(al_77f0ddfc[0]),
    .c(al_77f0ddfc[1]),
    .o(al_36605837));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_a6996a49 (
    .a(al_36605837),
    .b(al_643ac1f2),
    .c(al_68ba43d4),
    .o(al_39bb46f4));
  AL_MAP_LUT6 #(
    .EQN("(~E*~(~D*~B*~A*~(~F*C)))"),
    .INIT(64'h0000ffee0000fffe))
    al_c1a8b07b (
    .a(al_f80c5908),
    .b(al_39bb46f4),
    .c(al_12358921),
    .d(al_548d2e8d),
    .e(al_fdd1f60e),
    .f(al_af6614da),
    .o(al_17387d1));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*C*~B*A)"),
    .INIT(64'h0000000000000020))
    al_74afa4b (
    .a(al_1698ebe9),
    .b(al_85bba154),
    .c(al_6fa8f988),
    .d(al_20a6f635),
    .e(al_1d8c2b07),
    .f(al_56978088),
    .o(al_37f58acb));
  AL_MAP_LUT5 #(
    .EQN("(~(B)*~((~C*A))*~(D)*~(E)+B*~((~C*A))*~(D)*~(E)+B*~((~C*A))*D*~(E)+~(B)*~((~C*A))*~(D)*E+B*~((~C*A))*~(D)*E+B*(~C*A)*~(D)*E+B*~((~C*A))*D*E+B*(~C*A)*D*E)"),
    .INIT(32'hccfdc4f5))
    al_95c2e0d9 (
    .a(al_64e175a6),
    .b(al_bea385e7),
    .c(al_68ba43d4),
    .d(al_c925873),
    .e(al_21d722fe),
    .o(al_acb6d76c));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(D*C*~B))"),
    .INIT(16'hbaaa))
    al_9fda94f5 (
    .a(al_37f58acb),
    .b(al_acb6d76c),
    .c(al_8f22b7e0),
    .d(al_72403be8),
    .o(al_4421c6bd));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_6823225c (
    .a(al_c52cf3e8),
    .b(al_fdd1f60e),
    .o(al_1698ebe9));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_2fe9846b (
    .a(al_1698ebe9),
    .b(al_13f48428),
    .c(al_20a6f635),
    .d(al_cbafc250),
    .o(al_47b64b8f));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*B*~A)"),
    .INIT(32'h00000040))
    al_4b8dcf62 (
    .a(al_8afe6a9f),
    .b(al_72403be8),
    .c(al_ee3bb963),
    .d(al_548d2e8d),
    .e(al_cbafc250),
    .o(al_3c6cc34f));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~(A*~(D*C)))"),
    .INIT(16'hceee))
    al_b7b808db (
    .a(al_3c6cc34f),
    .b(al_47b64b8f),
    .c(al_907f6029),
    .d(al_d1e17be4),
    .o(al_4d7216c9));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    al_d4c341e7 (
    .a(al_20a6f635),
    .b(al_c52cf3e8),
    .c(al_1d8c2b07),
    .d(al_56978088),
    .o(al_1e340161));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(E*D*C*B))"),
    .INIT(32'heaaaaaaa))
    al_3645929c (
    .a(al_1e340161),
    .b(al_8f22b7e0),
    .c(al_6fa8f988),
    .d(al_13f48428),
    .e(al_c925873),
    .o(al_4be4ecdd));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*C*B*A)"),
    .INIT(32'h00008000))
    al_fdea729f (
    .a(al_8f22b7e0),
    .b(al_64e175a6),
    .c(al_6fa8f988),
    .d(al_13f48428),
    .e(al_c925873),
    .o(al_e04ba284));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_6c94f923 (
    .a(al_85bba154),
    .b(al_1d8c2b07),
    .c(al_56978088),
    .d(al_b348c1a2),
    .o(al_913e13a3));
  AL_MAP_LUT5 #(
    .EQN("(B*~(~D*~A*~(E*C)))"),
    .INIT(32'hccc8cc88))
    al_ba058319 (
    .a(al_e04ba284),
    .b(al_913e13a3),
    .c(al_20a6f635),
    .d(al_c52cf3e8),
    .e(al_bea385e7),
    .o(al_cf06a90));
  AL_MAP_LUT6 #(
    .EQN("(B*~(~(E*~D)*~(C*~(F*~A))))"),
    .INIT(64'h80cc8080c0ccc0c0))
    al_71d83145 (
    .a(al_8afe6a9f),
    .b(al_8f22b7e0),
    .c(al_64e175a6),
    .d(al_bea385e7),
    .e(al_c925873),
    .f(al_21d722fe),
    .o(al_4f19e5d0));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~(D*~B)*~(C*~A))"),
    .INIT(32'hffff7350))
    al_feace75b (
    .a(al_4f19e5d0),
    .b(al_85bba154),
    .c(al_13f48428),
    .d(al_fdd1f60e),
    .e(al_56978088),
    .o(al_da8b063f));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_e3736ab3 (
    .a(al_7fe117d0),
    .b(al_12358921),
    .o(al_531ee03c));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_502e5b0a (
    .a(al_177c7491),
    .b(al_5b769262),
    .o(al_4ba3ac36));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    al_be48396a (
    .a(al_531ee03c),
    .b(al_4ba3ac36),
    .c(al_72403be8),
    .d(al_fdd1f60e),
    .e(al_21d722fe),
    .o(al_92cc5462));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(E*~D)*~(~C*~B))"),
    .INIT(32'habffabab))
    al_d0ab896e (
    .a(al_f80c5908),
    .b(al_92cc5462),
    .c(al_2337d80f),
    .d(al_33f2071f),
    .e(al_e3f5d0d6),
    .o(al_3b1a77d7));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_8bd7a9ba (
    .a(al_2337d80f),
    .b(al_8f22b7e0),
    .o(al_4973ef09));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*~(B)*C*D*E)"),
    .INIT(32'h111105ff))
    al_fa910ae2 (
    .a(al_6fa8f988),
    .b(al_20a6f635),
    .c(al_c52cf3e8),
    .d(al_c35ead5c),
    .e(al_c925873),
    .o(al_638d20bb));
  AL_MAP_LUT6 #(
    .EQN("(B*~(~D*~(~C*~A*~(F*~E))))"),
    .INIT(64'hcc04cc00cc04cc04))
    al_6909d2ca (
    .a(al_638d20bb),
    .b(al_8f22b7e0),
    .c(al_64e175a6),
    .d(al_fdd1f60e),
    .e(al_bea385e7),
    .f(al_c925873),
    .o(al_b62e571a));
  AL_MAP_LUT6 #(
    .EQN("(~D*~(~F*~E*~C*B*~A))"),
    .INIT(64'h00ff00ff00ff00fb))
    al_584eb9d0 (
    .a(al_b62e571a),
    .b(al_d1e17be4),
    .c(al_edc29fee),
    .d(al_177c7491),
    .e(al_ea30f787),
    .f(al_cbafc250),
    .o(al_c59c6deb));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    al_9c845d60 (
    .a(al_24f8640d),
    .b(al_69f453c2),
    .c(al_cbafc250),
    .o(al_8f030415));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_18abf677 (
    .a(al_6b48ce98),
    .b(al_b984f6c1),
    .o(al_279c902b));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_e6bc7450 (
    .a(al_8afe6a9f),
    .b(al_85bba154),
    .c(al_fdd1f60e),
    .o(al_952d11ed));
  AL_MAP_LUT6 #(
    .EQN("(A*~(~F*~E*D*~C*~B))"),
    .INIT(64'haaaaaaaaaaaaa8aa))
    al_1b0e2519 (
    .a(al_952d11ed),
    .b(al_b156040b),
    .c(al_8aa33695),
    .d(al_51172105),
    .e(al_72403be8),
    .f(al_c52cf3e8),
    .o(al_24f8640d));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_b0c94024 (
    .a(al_a494216e),
    .b(al_fdd1f60e),
    .c(al_1d8c2b07),
    .d(al_56978088),
    .o(al_69f453c2));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    al_1a9fc9e1 (
    .a(al_24f8640d),
    .b(al_69f453c2),
    .c(al_3e886516),
    .d(al_e199650d),
    .o(al_6b2f12fa));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_9e0d9012 (
    .a(al_24ac8493[0]),
    .b(al_24ac8493[1]),
    .c(al_24ac8493[2]),
    .o(al_e1420a1f));
  AL_MAP_LUT6 #(
    .EQN("(~A*~(~E*~C*~(~F*~(~D*~B))))"),
    .INIT(64'h5555505055555554))
    al_1b7c1048 (
    .a(al_cbafc250),
    .b(al_e396ca5d),
    .c(al_48fcd383[2]),
    .d(al_e4dc5a7[1]),
    .e(al_f2f960a1),
    .f(al_c2463579),
    .o(al_8aa33695));
  AL_MAP_LUT6 #(
    .EQN("(~(~(F*D)*~(~E*B))*~(~C*~A))"),
    .INIT(64'hfa00fac80000c8c8))
    al_69da5d2d (
    .a(al_e1420a1f),
    .b(al_279c902b),
    .c(al_177c7491),
    .d(al_12358921),
    .e(al_cbafc250),
    .f(al_643ac1f2),
    .o(al_b156040b));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(~E*~D*~C*A))"),
    .INIT(32'h33333331))
    al_21453705 (
    .a(al_eb5c4882),
    .b(al_d75651de),
    .c(al_48fcd383[2]),
    .d(al_c925873),
    .e(al_f6643499),
    .o(al_51172105));
  AL_MAP_LUT4 #(
    .EQN("(~D*A*~(~C*~B))"),
    .INIT(16'h00a8))
    al_f369ac89 (
    .a(al_d1e17be4),
    .b(al_d27166fa),
    .c(al_6490a8fc),
    .d(al_48fcd383[1]),
    .o(al_8afe6a9f));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_5720f547 (
    .a(al_ee8473c1),
    .b(al_984d3b84[0]),
    .o(al_84a48183[0]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_7597f7be (
    .a(al_ee8473c1),
    .b(al_984d3b84[1]),
    .o(al_84a48183[1]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    al_eb1c8ede (
    .a(al_ee8473c1),
    .b(al_984d3b84[2]),
    .o(al_84a48183[2]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_d9a23bd2 (
    .a(al_ee8473c1),
    .b(al_984d3b84[3]),
    .o(al_84a48183[3]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    al_2162658d (
    .a(al_ee8473c1),
    .b(al_984d3b84[3]),
    .c(al_984d3b84[4]),
    .o(al_84a48183[4]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_347abbbd (
    .a(al_984d3b84[4]),
    .b(al_984d3b84[5]),
    .c(al_984d3b84[6]),
    .d(al_984d3b84[7]),
    .o(al_ab14fdf9));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~(~D*~C*~B)))"),
    .INIT(32'h0002aaaa))
    al_681307cf (
    .a(al_ab14fdf9),
    .b(al_984d3b84[0]),
    .c(al_984d3b84[1]),
    .d(al_984d3b84[2]),
    .e(al_984d3b84[3]),
    .o(al_25417591));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    al_46c13309 (
    .a(al_25417591),
    .b(al_d1e17be4),
    .c(al_d3482891),
    .o(al_ee8473c1));
  AL_MAP_LUT4 #(
    .EQN("(A*(D@(~C*~B)))"),
    .INIT(16'ha802))
    al_2d2fe367 (
    .a(al_ee8473c1),
    .b(al_984d3b84[3]),
    .c(al_984d3b84[4]),
    .d(al_984d3b84[5]),
    .o(al_84a48183[5]));
  AL_MAP_LUT5 #(
    .EQN("(A*(E@(~D*~C*~B)))"),
    .INIT(32'haaa80002))
    al_9ac2a76 (
    .a(al_ee8473c1),
    .b(al_984d3b84[3]),
    .c(al_984d3b84[4]),
    .d(al_984d3b84[5]),
    .e(al_984d3b84[6]),
    .o(al_84a48183[6]));
  AL_MAP_LUT6 #(
    .EQN("(F*A*~(~E*~D*~C*~B))"),
    .INIT(64'haaaaaaa800000000))
    al_3eebaff9 (
    .a(al_ee8473c1),
    .b(al_984d3b84[3]),
    .c(al_984d3b84[4]),
    .d(al_984d3b84[5]),
    .e(al_984d3b84[6]),
    .f(al_984d3b84[7]),
    .o(al_84a48183[7]));
  AL_MAP_LUT5 #(
    .EQN("(~D*A*~(~E*C*B))"),
    .INIT(32'h00aa002a))
    al_f20191e4 (
    .a(al_a1a0ec14),
    .b(al_2e2debcb),
    .c(al_cbafc250),
    .d(al_3e886516),
    .e(al_5f257019[5]),
    .o(al_a6c89001));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(E*~D*~C*~B))"),
    .INIT(32'haaabaaaa))
    al_8137a99f (
    .a(al_a6c89001),
    .b(al_85bba154),
    .c(al_a494216e),
    .d(al_fdd1f60e),
    .e(al_1d8c2b07),
    .o(al_81cdbd25));
  AL_MAP_LUT5 #(
    .EQN("~(B*~(~A*~(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)))"),
    .INIT(32'h33377377))
    al_7abe5540 (
    .a(al_907f6029),
    .b(al_d1e17be4),
    .c(al_edc29fee),
    .d(al_b1328a1f),
    .e(al_e5091a32),
    .o(al_ecd47e95));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_38d93521 (
    .a(al_b156040b),
    .b(al_51172105),
    .o(al_1f250659));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    al_679cc57 (
    .a(al_d1e17be4),
    .b(al_cbafc250),
    .c(al_1d8c2b07),
    .d(al_6490a8fc),
    .o(al_3557a617));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*~B)*~(D*~(~C*~A)))"),
    .INIT(32'hfb33fa00))
    al_622ad203 (
    .a(al_1f250659),
    .b(al_ecd47e95),
    .c(al_8aa33695),
    .d(al_3557a617),
    .e(al_d27166fa),
    .o(al_7ffb8465));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_39c52ca0 (
    .a(al_cbafc250),
    .b(al_f3f63e4d[0]),
    .o(al_630a3426[0]));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*C*~(B*A))"),
    .INIT(32'h00700000))
    al_e641b35d (
    .a(al_907f6029),
    .b(al_d1e17be4),
    .c(al_72403be8),
    .d(al_ee3bb963),
    .e(al_548d2e8d),
    .o(al_34d2745e));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(~E*~A*~(~C*B)))"),
    .INIT(32'h00ff00ae))
    al_54c9dbb7 (
    .a(al_f80c5908),
    .b(al_34d2745e),
    .c(al_ccc3c4e3),
    .d(al_fdd1f60e),
    .e(al_56978088),
    .o(al_e336c621));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_cc2776cc (
    .a(al_630a3426[0]),
    .b(al_f3f63e4d[1]),
    .o(al_a1a0ec14));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d1feb81 (
    .a(al_edc29fee),
    .b(al_3620963e),
    .c(al_1a7bad30),
    .o(al_907f6029));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_de90a103 (
    .a(al_5f257019[2]),
    .b(al_5f257019[3]),
    .c(al_5f257019[4]),
    .o(al_2e2debcb));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~D*~(~E*C*B)))"),
    .INIT(32'haa00aa80))
    al_c2aac481 (
    .a(al_a1a0ec14),
    .b(al_2e2debcb),
    .c(al_cbafc250),
    .d(al_3e886516),
    .e(al_5f257019[5]),
    .o(al_f80c5908));
  AL_MAP_LUT6 #(
    .EQN("(A*((D*~(E*C))*~(F)*~(B)+(D*~(E*C))*F*~(B)+~((D*~(E*C)))*F*B+(D*~(E*C))*F*B))"),
    .INIT(64'h8a88aa8802002200))
    al_1cd3f9a5 (
    .a(al_d1e17be4),
    .b(al_edc29fee),
    .c(al_1f6fed00),
    .d(al_b1328a1f),
    .e(al_beea368e),
    .f(al_e5091a32),
    .o(al_ccc3c4e3));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*~A)"),
    .INIT(8'hfe))
    al_e51cbd04 (
    .a(al_56978088),
    .b(al_6a534a0a),
    .c(al_4d3e0511),
    .o(al_b0eb70b2));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    al_fd79bf00 (
    .a(al_33f2071f),
    .b(al_24ac8493[0]),
    .o(al_63a836a9[0]));
  AL_MAP_LUT3 #(
    .EQN("~(A*(C@B))"),
    .INIT(8'hd7))
    al_a6dceeec (
    .a(al_33f2071f),
    .b(al_24ac8493[0]),
    .c(al_24ac8493[1]),
    .o(al_63a836a9[1]));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(D@(~C*~B)))"),
    .INIT(16'hfd57))
    al_a8f39433 (
    .a(al_33f2071f),
    .b(al_24ac8493[0]),
    .c(al_24ac8493[1]),
    .d(al_24ac8493[2]),
    .o(al_63a836a9[2]));
  AL_MAP_LUT6 #(
    .EQN("(A*~((D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))*~(E)*~(F)+A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)*~(E)*~(F)+A*~((D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))*E*~(F)+~(A)*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)*E*~(F)+A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)*E*~(F)+~(A)*~((D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))*~(E)*F+~(A)*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)*~(E)*F+~(A)*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)*E*F)"),
    .INIT(64'h51405555fbeaaaaa))
    al_84da321a (
    .a(al_5764731d),
    .b(al_d1e17be4),
    .c(al_edc29fee),
    .d(al_67d6ec64[0]),
    .e(al_33f2071f),
    .f(al_54d2aa3[0]),
    .o(al_c122424e[0]));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((~D*~B))*~(A)+C*(~D*~B)*~(A)+~(C)*(~D*~B)*A+C*(~D*~B)*A)"),
    .INIT(16'haf8d))
    al_e3504432 (
    .a(al_d1e17be4),
    .b(al_edc29fee),
    .c(al_67d6ec64[1]),
    .d(al_c925873),
    .o(al_dbee6318));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'hbf1510ba))
    al_33e63662 (
    .a(al_5764731d),
    .b(al_dbee6318),
    .c(al_33f2071f),
    .d(al_54d2aa3[0]),
    .e(al_54d2aa3[1]),
    .o(al_c122424e[1]));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~B))*~(A)+C*(D*~B)*~(A)+~(C)*(D*~B)*A+C*(D*~B)*A)"),
    .INIT(16'h8daf))
    al_a0145d13 (
    .a(al_d1e17be4),
    .b(al_edc29fee),
    .c(al_67d6ec64[2]),
    .d(al_c925873),
    .o(al_361cbc23));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~((~E*~D))*~(F)+A*~(B)*~(C)*(~E*~D)*~(F)+A*B*~(C)*(~E*~D)*~(F)+~(A)*~(B)*C*(~E*~D)*~(F)+A*~(B)*C*(~E*~D)*~(F)+A*B*C*(~E*~D)*~(F)+~(A)*~(B)*~(C)*~((~E*~D))*F+A*~(B)*~(C)*~((~E*~D))*F+~(A)*B*~(C)*~((~E*~D))*F+A*B*~(C)*~((~E*~D))*F+~(A)*~(B)*C*~((~E*~D))*F+A*~(B)*C*~((~E*~D))*F+A*B*C*~((~E*~D))*F+~(A)*~(B)*~(C)*(~E*~D)*F+~(A)*B*~(C)*(~E*~D)*F+~(A)*~(B)*C*(~E*~D)*F)"),
    .INIT(64'hbfbfbf15101010ba))
    al_d1dd248a (
    .a(al_5764731d),
    .b(al_361cbc23),
    .c(al_33f2071f),
    .d(al_54d2aa3[0]),
    .e(al_54d2aa3[1]),
    .f(al_54d2aa3[2]),
    .o(al_c122424e[2]));
  AL_MAP_LUT6 #(
    .EQN("(E*~((C*~((F*~B))*~(A)+C*(F*~B)*~(A)+~(C)*(F*~B)*A+C*(F*~B)*A))*~(D)+E*(C*~((F*~B))*~(A)+C*(F*~B)*~(A)+~(C)*(F*~B)*A+C*(F*~B)*A)*~(D)+~(E)*(C*~((F*~B))*~(A)+C*(F*~B)*~(A)+~(C)*(F*~B)*A+C*(F*~B)*A)*D+E*(C*~((F*~B))*~(A)+C*(F*~B)*~(A)+~(C)*(F*~B)*A+C*(F*~B)*A)*D)"),
    .INIT(64'h72ff720050ff5000))
    al_c411cc40 (
    .a(al_d1e17be4),
    .b(al_edc29fee),
    .c(al_67d6ec64[3]),
    .d(al_33f2071f),
    .e(al_54d2aa3[3]),
    .f(al_c925873),
    .o(al_6ec37834[3]));
  AL_MAP_LUT6 #(
    .EQN("(B*~((F@(~E*~D*~C)))*~(A)+B*(F@(~E*~D*~C))*~(A)+~(B)*(F@(~E*~D*~C))*A+B*(F@(~E*~D*~C))*A)"),
    .INIT(64'heeeeeee44444444e))
    al_67419235 (
    .a(al_5764731d),
    .b(al_6ec37834[3]),
    .c(al_54d2aa3[0]),
    .d(al_54d2aa3[1]),
    .e(al_54d2aa3[2]),
    .f(al_54d2aa3[3]),
    .o(al_c122424e[3]));
  AL_MAP_LUT6 #(
    .EQN("(A*B*~((D*~C))*~(E)*~(F)+A*B*(D*~C)*~(E)*~(F)+A*B*~((D*~C))*E*~(F)+~(A)*~(B)*(D*~C)*E*~(F)+~(A)*B*(D*~C)*E*~(F)+A*B*(D*~C)*E*~(F)+~(A)*~(B)*~((D*~C))*~(E)*F+A*~(B)*~((D*~C))*~(E)*F+~(A)*B*~((D*~C))*~(E)*F+~(A)*~(B)*(D*~C)*~(E)*F+A*~(B)*(D*~C)*~(E)*F+~(A)*B*(D*~C)*~(E)*F+A*~(B)*~((D*~C))*E*F+~(A)*~(B)*(D*~C)*E*F+A*~(B)*(D*~C)*E*F+~(A)*B*(D*~C)*E*F)"),
    .INIT(64'h272277778d888888))
    al_6d30852c (
    .a(al_5764731d),
    .b(al_d10bb6dd),
    .c(al_d1e17be4),
    .d(al_67d6ec64[4]),
    .e(al_33f2071f),
    .f(al_54d2aa3[4]),
    .o(al_c122424e[4]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_8d4c3e2f (
    .a(al_54d2aa3[0]),
    .b(al_54d2aa3[1]),
    .c(al_54d2aa3[2]),
    .d(al_54d2aa3[3]),
    .o(al_d10bb6dd));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_7c4f6716 (
    .a(al_d10bb6dd),
    .b(al_54d2aa3[4]),
    .o(al_95e117eb));
  AL_MAP_LUT6 #(
    .EQN("(A*B*~((D*~C))*~(E)*~(F)+A*B*(D*~C)*~(E)*~(F)+A*B*~((D*~C))*E*~(F)+~(A)*~(B)*(D*~C)*E*~(F)+~(A)*B*(D*~C)*E*~(F)+A*B*(D*~C)*E*~(F)+~(A)*~(B)*~((D*~C))*~(E)*F+A*~(B)*~((D*~C))*~(E)*F+~(A)*B*~((D*~C))*~(E)*F+~(A)*~(B)*(D*~C)*~(E)*F+A*~(B)*(D*~C)*~(E)*F+~(A)*B*(D*~C)*~(E)*F+A*~(B)*~((D*~C))*E*F+~(A)*~(B)*(D*~C)*E*F+A*~(B)*(D*~C)*E*F+~(A)*B*(D*~C)*E*F)"),
    .INIT(64'h272277778d888888))
    al_6fc8817d (
    .a(al_5764731d),
    .b(al_95e117eb),
    .c(al_d1e17be4),
    .d(al_67d6ec64[5]),
    .e(al_33f2071f),
    .f(al_54d2aa3[5]),
    .o(al_c122424e[5]));
  AL_MAP_LUT6 #(
    .EQN("(A*B*~((D*~C))*~(E)*~(F)+A*B*(D*~C)*~(E)*~(F)+A*B*~((D*~C))*E*~(F)+~(A)*~(B)*(D*~C)*E*~(F)+~(A)*B*(D*~C)*E*~(F)+A*B*(D*~C)*E*~(F)+~(A)*~(B)*~((D*~C))*~(E)*F+A*~(B)*~((D*~C))*~(E)*F+~(A)*B*~((D*~C))*~(E)*F+~(A)*~(B)*(D*~C)*~(E)*F+A*~(B)*(D*~C)*~(E)*F+~(A)*B*(D*~C)*~(E)*F+A*~(B)*~((D*~C))*E*F+~(A)*~(B)*(D*~C)*E*F+A*~(B)*(D*~C)*E*F+~(A)*B*(D*~C)*E*F)"),
    .INIT(64'h272277778d888888))
    al_57e451a5 (
    .a(al_5764731d),
    .b(al_eeaafdd6),
    .c(al_d1e17be4),
    .d(al_67d6ec64[6]),
    .e(al_33f2071f),
    .f(al_54d2aa3[6]),
    .o(al_c122424e[6]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_50bf4e22 (
    .a(al_54d2aa3[0]),
    .b(al_54d2aa3[1]),
    .c(al_54d2aa3[2]),
    .d(al_54d2aa3[3]),
    .e(al_54d2aa3[4]),
    .f(al_54d2aa3[5]),
    .o(al_eeaafdd6));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_223d8913 (
    .a(al_eeaafdd6),
    .b(al_54d2aa3[6]),
    .o(al_af3a6b91));
  AL_MAP_LUT5 #(
    .EQN("(~D*~C*~B*~(~E*A))"),
    .INIT(32'h00030001))
    al_4672f984 (
    .a(al_af3a6b91),
    .b(al_1698ebe9),
    .c(al_56978088),
    .d(al_c388f857),
    .e(al_54d2aa3[7]),
    .o(al_5764731d));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*(D*~C)*E*~(F)+~(A)*B*(D*~C)*E*~(F)+~(A)*~(B)*~((D*~C))*~(E)*F+A*~(B)*~((D*~C))*~(E)*F+~(A)*B*~((D*~C))*~(E)*F+~(A)*~(B)*(D*~C)*~(E)*F+A*~(B)*(D*~C)*~(E)*F+~(A)*B*(D*~C)*~(E)*F+A*~(B)*~((D*~C))*E*F+~(A)*~(B)*(D*~C)*E*F+A*~(B)*(D*~C)*E*F+~(A)*B*(D*~C)*E*F)"),
    .INIT(64'h2722777705000000))
    al_d9782e47 (
    .a(al_5764731d),
    .b(al_af3a6b91),
    .c(al_d1e17be4),
    .d(al_67d6ec64[7]),
    .e(al_33f2071f),
    .f(al_54d2aa3[7]),
    .o(al_c122424e[7]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_bebac684 (
    .a(al_af3a6b91),
    .b(al_fdd1f60e),
    .c(al_54d2aa3[7]),
    .o(al_114ce5a4));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    al_4de7da09 (
    .a(al_5b769262),
    .b(al_77f0ddfc[0]),
    .o(al_b3968bab[0]));
  AL_MAP_LUT3 #(
    .EQN("~(A*(C@B))"),
    .INIT(8'hd7))
    al_cef218ce (
    .a(al_5b769262),
    .b(al_77f0ddfc[0]),
    .c(al_77f0ddfc[1]),
    .o(al_b3968bab[1]));
  AL_MAP_LUT3 #(
    .EQN("~(A*(C@B))"),
    .INIT(8'hd7))
    al_edacd113 (
    .a(al_cbafc250),
    .b(al_f3f63e4d[0]),
    .c(al_f3f63e4d[1]),
    .o(al_630a3426[1]));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT(16'hddf5))
    al_4811759a (
    .a(al_1d8c2b07),
    .b(al_e8bb9040[0]),
    .c(al_acbf9207[0]),
    .d(al_4fb6999c),
    .o(al_77695f5b[0]));
  AL_MAP_LUT6 #(
    .EQN("~((F*A*~(E*D))*~(C)*~(B)+(F*A*~(E*D))*C*~(B)+~((F*A*~(E*D)))*C*B+(F*A*~(E*D))*C*B)"),
    .INIT(64'h3f1d1d1d3f3f3f3f))
    al_a2155a16 (
    .a(al_edc29fee),
    .b(al_1d8c2b07),
    .c(al_e8bb9040[10]),
    .d(al_5f257019[4]),
    .e(al_5f257019[5]),
    .f(al_6c9db937[4]),
    .o(al_bb4cafc));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~((~C*B))*~(D)*~(E)*~(F)+~(A)*(~C*B)*~(D)*~(E)*~(F)+A*(~C*B)*~(D)*~(E)*~(F)+~(A)*~((~C*B))*~(D)*E*~(F)+~(A)*(~C*B)*~(D)*E*~(F)+A*(~C*B)*~(D)*E*~(F)+~(A)*~((~C*B))*D*E*~(F)+A*~((~C*B))*D*E*~(F)+~(A)*(~C*B)*D*E*~(F)+A*(~C*B)*D*E*~(F)+~(A)*~((~C*B))*~(D)*~(E)*F+~(A)*(~C*B)*~(D)*~(E)*F+A*(~C*B)*~(D)*~(E)*F+~(A)*~((~C*B))*D*~(E)*F+~(A)*(~C*B)*D*~(E)*F+~(A)*~((~C*B))*~(D)*E*F+~(A)*(~C*B)*~(D)*E*F+A*(~C*B)*~(D)*E*F+~(A)*~((~C*B))*D*E*F+~(A)*(~C*B)*D*E*F)"),
    .INIT(64'h555d555dff5d005d))
    al_da15a503 (
    .a(al_bb4cafc),
    .b(al_6e9a1ae[1]),
    .c(al_edc29fee),
    .d(al_1d8c2b07),
    .e(al_acbf9207[10]),
    .f(al_4fb6999c),
    .o(al_77695f5b[10]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*A))"),
    .INIT(16'h7f00))
    al_303b0074 (
    .a(al_5f257019[3]),
    .b(al_5f257019[4]),
    .c(al_5f257019[5]),
    .d(al_6c9db937[2]),
    .o(al_6e9a1ae[2]));
  AL_MAP_LUT5 #(
    .EQN("(E*~(D*~(~C*~(B*A))))"),
    .INIT(32'h07ff0000))
    al_1565140e (
    .a(al_5f257019[2]),
    .b(al_5f257019[3]),
    .c(al_5f257019[4]),
    .d(al_5f257019[5]),
    .e(al_6c9db937[5]),
    .o(al_6e9a1ae[5]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    al_dc89cd3e (
    .a(al_6e9a1ae[5]),
    .b(al_6e9a1ae[2]),
    .c(al_edc29fee),
    .o(al_4f97dd8c));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((D*~(C)*~(E)+D*C*~(E)+~(D)*C*E+D*C*E))*~(B)+~A*(D*~(C)*~(E)+D*C*~(E)+~(D)*C*E+D*C*E)*~(B)+~(~A)*(D*~(C)*~(E)+D*C*~(E)+~(D)*C*E+D*C*E)*B+~A*(D*~(C)*~(E)+D*C*~(E)+~(D)*C*E+D*C*E)*B)"),
    .INIT(32'hd1d1dd11))
    al_4a63ff33 (
    .a(al_4f97dd8c),
    .b(al_1d8c2b07),
    .c(al_e8bb9040[11]),
    .d(al_acbf9207[11]),
    .e(al_4fb6999c),
    .o(al_77695f5b[11]));
  AL_MAP_LUT4 #(
    .EQN("~(A*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT(16'h775f))
    al_1d9e0733 (
    .a(al_1d8c2b07),
    .b(al_e8bb9040[12]),
    .c(al_acbf9207[12]),
    .d(al_4fb6999c),
    .o(al_d0ab12fe));
  AL_MAP_LUT5 #(
    .EQN("~(C*~(~E*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    .INIT(32'h0f0fcfaf))
    al_a9a7588c (
    .a(al_6e9a1ae[3]),
    .b(al_6e9a1ae[6]),
    .c(al_d0ab12fe),
    .d(al_edc29fee),
    .e(al_1d8c2b07),
    .o(al_77695f5b[12]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*~A))"),
    .INIT(8'hb0))
    al_5484a280 (
    .a(al_2e2debcb),
    .b(al_5f257019[5]),
    .c(al_6c9db937[7]),
    .o(al_6e9a1ae[7]));
  AL_MAP_LUT6 #(
    .EQN("~((F*~A*~(E*D))*~(C)*~(B)+(F*~A*~(E*D))*C*~(B)+~((F*~A*~(E*D)))*C*B+(F*~A*~(E*D))*C*B)"),
    .INIT(64'h3f2e2e2e3f3f3f3f))
    al_1eabfaac (
    .a(al_edc29fee),
    .b(al_1d8c2b07),
    .c(al_e8bb9040[13]),
    .d(al_5f257019[4]),
    .e(al_5f257019[5]),
    .f(al_6c9db937[4]),
    .o(al_a48c9e07));
  AL_MAP_LUT6 #(
    .EQN("(~(B)*~((C*A))*~(D)*~(E)*~(F)+~(B)*(C*A)*~(D)*~(E)*~(F)+B*(C*A)*~(D)*~(E)*~(F)+~(B)*~((C*A))*~(D)*E*~(F)+~(B)*(C*A)*~(D)*E*~(F)+B*(C*A)*~(D)*E*~(F)+~(B)*~((C*A))*D*E*~(F)+B*~((C*A))*D*E*~(F)+~(B)*(C*A)*D*E*~(F)+B*(C*A)*D*E*~(F)+~(B)*~((C*A))*~(D)*~(E)*F+~(B)*(C*A)*~(D)*~(E)*F+B*(C*A)*~(D)*~(E)*F+~(B)*~((C*A))*D*~(E)*F+~(B)*(C*A)*D*~(E)*F+~(B)*~((C*A))*~(D)*E*F+~(B)*(C*A)*~(D)*E*F+B*(C*A)*~(D)*E*F+~(B)*~((C*A))*D*E*F+~(B)*(C*A)*D*E*F)"),
    .INIT(64'h33b333b3ffb300b3))
    al_75b4abc7 (
    .a(al_6e9a1ae[7]),
    .b(al_a48c9e07),
    .c(al_edc29fee),
    .d(al_1d8c2b07),
    .e(al_acbf9207[13]),
    .f(al_4fb6999c),
    .o(al_77695f5b[13]));
  AL_MAP_LUT4 #(
    .EQN("~(A*~((D*~C))*~(B)+A*(D*~C)*~(B)+~(A)*(D*~C)*B+A*(D*~C)*B)"),
    .INIT(16'hd1dd))
    al_ae603fe7 (
    .a(al_6e9a1ae[5]),
    .b(al_edc29fee),
    .c(al_5f257019[5]),
    .d(al_6c9db937[8]),
    .o(al_88a372db));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((D*~(C)*~(E)+D*C*~(E)+~(D)*C*E+D*C*E))*~(B)+~A*(D*~(C)*~(E)+D*C*~(E)+~(D)*C*E+D*C*E)*~(B)+~(~A)*(D*~(C)*~(E)+D*C*~(E)+~(D)*C*E+D*C*E)*B+~A*(D*~(C)*~(E)+D*C*~(E)+~(D)*C*E+D*C*E)*B)"),
    .INIT(32'hd1d1dd11))
    al_f8a4925f (
    .a(al_88a372db),
    .b(al_1d8c2b07),
    .c(al_e8bb9040[14]),
    .d(al_acbf9207[14]),
    .e(al_4fb6999c),
    .o(al_77695f5b[14]));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~(C*B*A))"),
    .INIT(32'h007f0000))
    al_9422667f (
    .a(al_5f257019[2]),
    .b(al_5f257019[3]),
    .c(al_5f257019[4]),
    .d(al_5f257019[5]),
    .e(al_6c9db937[9]),
    .o(al_6e9a1ae[9]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~(~B*~A)))"),
    .INIT(16'h1f00))
    al_e28a9a76 (
    .a(al_5f257019[3]),
    .b(al_5f257019[4]),
    .c(al_5f257019[5]),
    .d(al_6c9db937[6]),
    .o(al_6e9a1ae[6]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    al_2de3b749 (
    .a(al_6e9a1ae[9]),
    .b(al_6e9a1ae[6]),
    .c(al_edc29fee),
    .o(al_fbb2ea7a));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((D*~(C)*~(E)+D*C*~(E)+~(D)*C*E+D*C*E))*~(B)+~A*(D*~(C)*~(E)+D*C*~(E)+~(D)*C*E+D*C*E)*~(B)+~(~A)*(D*~(C)*~(E)+D*C*~(E)+~(D)*C*E+D*C*E)*B+~A*(D*~(C)*~(E)+D*C*~(E)+~(D)*C*E+D*C*E)*B)"),
    .INIT(32'hd1d1dd11))
    al_439c9ff1 (
    .a(al_fbb2ea7a),
    .b(al_1d8c2b07),
    .c(al_e8bb9040[15]),
    .d(al_acbf9207[15]),
    .e(al_4fb6999c),
    .o(al_77695f5b[15]));
  AL_MAP_LUT6 #(
    .EQN("((~B*A)*~((E*~(D)*~(F)+E*D*~(F)+~(E)*D*F+E*D*F))*~(C)+(~B*A)*(E*~(D)*~(F)+E*D*~(F)+~(E)*D*F+E*D*F)*~(C)+~((~B*A))*(E*~(D)*~(F)+E*D*~(F)+~(E)*D*F+E*D*F)*C+(~B*A)*(E*~(D)*~(F)+E*D*~(F)+~(E)*D*F+E*D*F)*C)"),
    .INIT(64'hf202f202f2f20202))
    al_f2588bcf (
    .a(al_6e9a1ae[7]),
    .b(al_edc29fee),
    .c(al_1d8c2b07),
    .d(al_e8bb9040[16]),
    .e(al_acbf9207[16]),
    .f(al_4fb6999c),
    .o(al_77695f5b[16]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    al_781702a3 (
    .a(al_e8bb9040[17]),
    .b(al_acbf9207[17]),
    .c(al_4fb6999c),
    .o(al_36d5f4c5));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*~D*~B)*~(A)*~(C)+~(E*~D*~B)*A*~(C)+~(~(E*~D*~B))*A*C+~(E*~D*~B)*A*C)"),
    .INIT(32'h50535050))
    al_4d5c3cd4 (
    .a(al_36d5f4c5),
    .b(al_edc29fee),
    .c(al_1d8c2b07),
    .d(al_5f257019[5]),
    .e(al_6c9db937[8]),
    .o(al_77695f5b[17]));
  AL_MAP_LUT6 #(
    .EQN("((~B*A)*~((E*~(D)*~(F)+E*D*~(F)+~(E)*D*F+E*D*F))*~(C)+(~B*A)*(E*~(D)*~(F)+E*D*~(F)+~(E)*D*F+E*D*F)*~(C)+~((~B*A))*(E*~(D)*~(F)+E*D*~(F)+~(E)*D*F+E*D*F)*C+(~B*A)*(E*~(D)*~(F)+E*D*~(F)+~(E)*D*F+E*D*F)*C)"),
    .INIT(64'hf202f202f2f20202))
    al_e7ec6efc (
    .a(al_6e9a1ae[9]),
    .b(al_edc29fee),
    .c(al_1d8c2b07),
    .d(al_e8bb9040[18]),
    .e(al_acbf9207[18]),
    .f(al_4fb6999c),
    .o(al_77695f5b[18]));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT(16'hddf5))
    al_dbee17e5 (
    .a(al_1d8c2b07),
    .b(al_e8bb9040[1]),
    .c(al_acbf9207[1]),
    .d(al_4fb6999c),
    .o(al_77695f5b[1]));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT(16'hddf5))
    al_afec4398 (
    .a(al_1d8c2b07),
    .b(al_e8bb9040[2]),
    .c(al_acbf9207[2]),
    .d(al_4fb6999c),
    .o(al_77695f5b[2]));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT(16'hddf5))
    al_97e0040b (
    .a(al_1d8c2b07),
    .b(al_e8bb9040[3]),
    .c(al_acbf9207[3]),
    .d(al_4fb6999c),
    .o(al_77695f5b[3]));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT(16'hddf5))
    al_364e4091 (
    .a(al_1d8c2b07),
    .b(al_e8bb9040[4]),
    .c(al_acbf9207[4]),
    .d(al_4fb6999c),
    .o(al_77695f5b[4]));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT(16'hddf5))
    al_d0f9845f (
    .a(al_1d8c2b07),
    .b(al_e8bb9040[5]),
    .c(al_acbf9207[5]),
    .d(al_4fb6999c),
    .o(al_77695f5b[5]));
  AL_MAP_LUT6 #(
    .EQN("(~(~F*A)*~((D*~(C)*~(E)+D*C*~(E)+~(D)*C*E+D*C*E))*~(B)+~(~F*A)*(D*~(C)*~(E)+D*C*~(E)+~(D)*C*E+D*C*E)*~(B)+~(~(~F*A))*(D*~(C)*~(E)+D*C*~(E)+~(D)*C*E+D*C*E)*B+~(~F*A)*(D*~(C)*~(E)+D*C*~(E)+~(D)*C*E+D*C*E)*B)"),
    .INIT(64'hf3f3ff33d1d1dd11))
    al_4579afb5 (
    .a(al_edc29fee),
    .b(al_1d8c2b07),
    .c(al_e8bb9040[6]),
    .d(al_acbf9207[6]),
    .e(al_4fb6999c),
    .f(al_6c9db937[0]),
    .o(al_77695f5b[6]));
  AL_MAP_LUT5 #(
    .EQN("(E*~(D*C*B*A))"),
    .INIT(32'h7fff0000))
    al_7f66479d (
    .a(al_5f257019[2]),
    .b(al_5f257019[3]),
    .c(al_5f257019[4]),
    .d(al_5f257019[5]),
    .e(al_6c9db937[1]),
    .o(al_6e9a1ae[1]));
  AL_MAP_LUT6 #(
    .EQN("(~(B*~A)*~((E*~(D)*~(F)+E*D*~(F)+~(E)*D*F+E*D*F))*~(C)+~(B*~A)*(E*~(D)*~(F)+E*D*~(F)+~(E)*D*F+E*D*F)*~(C)+~(~(B*~A))*(E*~(D)*~(F)+E*D*~(F)+~(E)*D*F+E*D*F)*C+~(B*~A)*(E*~(D)*~(F)+E*D*~(F)+~(E)*D*F+E*D*F)*C)"),
    .INIT(64'hfb0bfb0bfbfb0b0b))
    al_8e61b8d8 (
    .a(al_6e9a1ae[1]),
    .b(al_edc29fee),
    .c(al_1d8c2b07),
    .d(al_e8bb9040[7]),
    .e(al_acbf9207[7]),
    .f(al_4fb6999c),
    .o(al_77695f5b[7]));
  AL_MAP_LUT6 #(
    .EQN("(~(B*~A)*~((E*~(D)*~(F)+E*D*~(F)+~(E)*D*F+E*D*F))*~(C)+~(B*~A)*(E*~(D)*~(F)+E*D*~(F)+~(E)*D*F+E*D*F)*~(C)+~(~(B*~A))*(E*~(D)*~(F)+E*D*~(F)+~(E)*D*F+E*D*F)*C+~(B*~A)*(E*~(D)*~(F)+E*D*~(F)+~(E)*D*F+E*D*F)*C)"),
    .INIT(64'hfb0bfb0bfbfb0b0b))
    al_b1220d55 (
    .a(al_6e9a1ae[2]),
    .b(al_edc29fee),
    .c(al_1d8c2b07),
    .d(al_e8bb9040[8]),
    .e(al_acbf9207[8]),
    .f(al_4fb6999c),
    .o(al_77695f5b[8]));
  AL_MAP_LUT5 #(
    .EQN("(E*~(D*C*~(~B*~A)))"),
    .INIT(32'h1fff0000))
    al_72a91bf7 (
    .a(al_5f257019[2]),
    .b(al_5f257019[3]),
    .c(al_5f257019[4]),
    .d(al_5f257019[5]),
    .e(al_6c9db937[3]),
    .o(al_6e9a1ae[3]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    al_ad750a8c (
    .a(al_6e9a1ae[3]),
    .b(al_edc29fee),
    .c(al_6c9db937[0]),
    .o(al_9dbb5412));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((D*~(C)*~(E)+D*C*~(E)+~(D)*C*E+D*C*E))*~(B)+~A*(D*~(C)*~(E)+D*C*~(E)+~(D)*C*E+D*C*E)*~(B)+~(~A)*(D*~(C)*~(E)+D*C*~(E)+~(D)*C*E+D*C*E)*B+~A*(D*~(C)*~(E)+D*C*~(E)+~(D)*C*E+D*C*E)*B)"),
    .INIT(32'hd1d1dd11))
    al_99be4668 (
    .a(al_9dbb5412),
    .b(al_1d8c2b07),
    .c(al_e8bb9040[9]),
    .d(al_acbf9207[9]),
    .e(al_4fb6999c),
    .o(al_77695f5b[9]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(D@(~C*B)))"),
    .INIT(16'hfbae))
    al_470bcfd9 (
    .a(al_8e6b9688),
    .b(al_cbafc250),
    .c(al_3e886516),
    .d(al_5f257019[0]),
    .o(al_20b55994[0]));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(E@(~D*~C*B)))"),
    .INIT(32'hfffbaaae))
    al_142b5f69 (
    .a(al_8e6b9688),
    .b(al_cbafc250),
    .c(al_3e886516),
    .d(al_5f257019[0]),
    .e(al_5f257019[1]),
    .o(al_20b55994[1]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+~(A)*B*~(C)+A*B*~(C)+~(A)*~(B)*C+A*~(B)*C)"),
    .INIT(8'h3e))
    al_911ffca9 (
    .a(al_8e6b9688),
    .b(al_aa5dc84f),
    .c(al_5f257019[2]),
    .o(al_20b55994[2]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(D@(~C*B)))"),
    .INIT(16'hfbae))
    al_c6f47203 (
    .a(al_8e6b9688),
    .b(al_aa5dc84f),
    .c(al_5f257019[2]),
    .d(al_5f257019[3]),
    .o(al_20b55994[3]));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(E@(~D*~C*B)))"),
    .INIT(32'hfffbaaae))
    al_e4f22c90 (
    .a(al_8e6b9688),
    .b(al_aa5dc84f),
    .c(al_5f257019[2]),
    .d(al_5f257019[3]),
    .e(al_5f257019[4]),
    .o(al_20b55994[4]));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*~A))"),
    .INIT(16'hf3a2))
    al_32e38c55 (
    .a(al_85bba154),
    .b(al_cbafc250),
    .c(al_3e886516),
    .d(al_f28e4921),
    .o(al_8e6b9688));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    al_9157d647 (
    .a(al_cbafc250),
    .b(al_3e886516),
    .c(al_5f257019[0]),
    .d(al_5f257019[1]),
    .o(al_aa5dc84f));
  AL_MAP_LUT4 #(
    .EQN("(A*~((C*B))*~(D)+~(A)*(C*B)*~(D)+A*(C*B)*~(D)+~(A)*~((C*B))*D+A*~((C*B))*D)"),
    .INIT(16'h3fea))
    al_f465ea04 (
    .a(al_8e6b9688),
    .b(al_aa5dc84f),
    .c(al_2e2debcb),
    .d(al_5f257019[5]),
    .o(al_20b55994[5]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .INIT(16'h4540))
    al_b2d117 (
    .a(al_a12adb97),
    .b(al_e512aff[0]),
    .c(al_e512aff[14]),
    .d(al_f5f472e[0]),
    .o(al_c007c6a1[0]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .INIT(16'h4540))
    al_d8ee22eb (
    .a(al_a12adb97),
    .b(al_e512aff[10]),
    .c(al_e512aff[14]),
    .d(al_f5f472e[10]),
    .o(al_c007c6a1[10]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .INIT(16'h4540))
    al_3fcf77a4 (
    .a(al_a12adb97),
    .b(al_e512aff[11]),
    .c(al_e512aff[14]),
    .d(al_f5f472e[11]),
    .o(al_c007c6a1[11]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .INIT(16'h4540))
    al_ee5824fa (
    .a(al_a12adb97),
    .b(al_e512aff[12]),
    .c(al_e512aff[14]),
    .d(al_f5f472e[12]),
    .o(al_c007c6a1[12]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    al_d7bac4fb (
    .a(al_4ba3ac36),
    .b(al_7fe117d0),
    .c(al_6fa8f988),
    .d(al_20a6f635),
    .o(al_a12adb97));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .INIT(16'h4540))
    al_a86f7fe (
    .a(al_a12adb97),
    .b(al_e512aff[13]),
    .c(al_e512aff[14]),
    .d(al_f5f472e[13]),
    .o(al_c007c6a1[13]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    al_f6f8bb46 (
    .a(al_a12adb97),
    .b(al_e512aff[14]),
    .c(al_f5f472e[14]),
    .o(al_c007c6a1[14]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .INIT(16'h4540))
    al_82655128 (
    .a(al_a12adb97),
    .b(al_e512aff[1]),
    .c(al_e512aff[14]),
    .d(al_f5f472e[1]),
    .o(al_c007c6a1[1]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)*~(E)*~(A)+(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)*E*~(A)+~((D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))*E*A+(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)*E*A)"),
    .INIT(32'hefea4540))
    al_cbe2a894 (
    .a(al_a12adb97),
    .b(al_e512aff[2]),
    .c(al_e512aff[14]),
    .d(al_f5f472e[2]),
    .e(al_af6614da),
    .o(al_c007c6a1[2]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .INIT(16'h4540))
    al_19a600da (
    .a(al_a12adb97),
    .b(al_e512aff[3]),
    .c(al_e512aff[14]),
    .d(al_f5f472e[3]),
    .o(al_c007c6a1[3]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .INIT(16'h4540))
    al_36d3e2f5 (
    .a(al_a12adb97),
    .b(al_e512aff[4]),
    .c(al_e512aff[14]),
    .d(al_f5f472e[4]),
    .o(al_c007c6a1[4]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .INIT(16'h4540))
    al_604a2be6 (
    .a(al_a12adb97),
    .b(al_e512aff[5]),
    .c(al_e512aff[14]),
    .d(al_f5f472e[5]),
    .o(al_c007c6a1[5]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .INIT(16'h4540))
    al_8072918 (
    .a(al_a12adb97),
    .b(al_e512aff[6]),
    .c(al_e512aff[14]),
    .d(al_f5f472e[6]),
    .o(al_c007c6a1[6]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .INIT(16'h4540))
    al_7fd0a175 (
    .a(al_a12adb97),
    .b(al_e512aff[7]),
    .c(al_e512aff[14]),
    .d(al_f5f472e[7]),
    .o(al_c007c6a1[7]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .INIT(16'h4540))
    al_d61e0086 (
    .a(al_a12adb97),
    .b(al_e512aff[8]),
    .c(al_e512aff[14]),
    .d(al_f5f472e[8]),
    .o(al_c007c6a1[8]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .INIT(16'h4540))
    al_2443d423 (
    .a(al_a12adb97),
    .b(al_e512aff[9]),
    .c(al_e512aff[14]),
    .d(al_f5f472e[9]),
    .o(al_c007c6a1[9]));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*~B)*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(32'hf7b3f5a0))
    al_5305f2a7 (
    .a(al_edc29fee),
    .b(al_33f2071f),
    .c(al_e512aff[6]),
    .d(al_e512aff[9]),
    .e(al_bea385e7),
    .o(al_4a89f542));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*~A))"),
    .INIT(8'hdc))
    al_71ccec (
    .a(al_33f2071f),
    .b(al_e512aff[6]),
    .c(al_642e830e),
    .o(al_70a59d2e));
  AL_MAP_LUT5 #(
    .EQN("(~(E@C)*(~(A)*~(B)*~(D)+A*B*D))"),
    .INIT(32'h80100801))
    al_c6d9a076 (
    .a(al_e512aff[2]),
    .b(al_e512aff[3]),
    .c(al_e512aff[4]),
    .d(al_19bf88c2[2]),
    .e(al_19bf88c2[4]),
    .o(al_a8d1cf64));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*~B*~A)"),
    .INIT(64'h1000000000000000))
    al_66ff6e9b (
    .a(al_fdd1f60e),
    .b(al_e512aff[0]),
    .c(al_e512aff[1]),
    .d(al_e512aff[5]),
    .e(al_e512aff[6]),
    .f(al_e512aff[7]),
    .o(al_1751a6d0));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    al_f2e7663f (
    .a(al_e512aff[8]),
    .b(al_e512aff[9]),
    .c(al_e512aff[10]),
    .d(al_e512aff[11]),
    .o(al_360cb20));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*C*B*A)"),
    .INIT(64'h0000000000000080))
    al_e1a3c1b6 (
    .a(al_1751a6d0),
    .b(al_a8d1cf64),
    .c(al_360cb20),
    .d(al_e512aff[12]),
    .e(al_e512aff[13]),
    .f(al_e512aff[14]),
    .o(al_eaacfd93));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(~A*~(E*~(D*~B))))"),
    .INIT(32'h0e0f0a0a))
    al_b90b89c3 (
    .a(al_eaacfd93),
    .b(al_1698ebe9),
    .c(al_ea441981),
    .d(al_c35ead5c),
    .e(al_643ac1f2),
    .o(al_ffd3f5d1));
  AL_MAP_LUT6 #(
    .EQN("(F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000100000000))
    al_b3fbe1a6 (
    .a(al_bff87853[1]),
    .b(al_bff87853[2]),
    .c(al_bff87853[4]),
    .d(al_bff87853[5]),
    .e(al_bff87853[6]),
    .f(al_bff87853[7]),
    .o(al_96d069e8));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_c1604fa0 (
    .a(al_bff87853[8]),
    .b(al_bff87853[9]),
    .c(al_bff87853[10]),
    .d(al_bff87853[12]),
    .o(al_68e39bd9));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    al_fe6e504e (
    .a(al_96d069e8),
    .b(al_68e39bd9),
    .c(al_bff87853[13]),
    .d(al_bff87853[14]),
    .e(al_bff87853[15]),
    .o(al_a140f198));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*B*A)"),
    .INIT(32'h00000080))
    al_b5fb917d (
    .a(al_a140f198),
    .b(al_f731da11),
    .c(al_bff87853[0]),
    .d(al_bff87853[3]),
    .e(al_bff87853[11]),
    .o(al_d09ba8fa));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    al_54dae24d (
    .a(al_d09ba8fa),
    .o(al_ae339d26[2]));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D*~B*~A))"),
    .INIT(16'hf1f0))
    al_ea57c117 (
    .a(al_85bba154),
    .b(al_33f2071f),
    .c(al_12358921),
    .d(al_68ba43d4),
    .o(al_4fe9a477));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    al_cf24ad56 (
    .a(al_d1e17be4),
    .b(al_edc29fee),
    .c(al_beea368e),
    .o(al_8f22b7e0));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_f61ea9c6 (
    .a(al_821706b3[4]),
    .b(al_821706b3[5]),
    .c(al_821706b3[7]),
    .d(al_821706b3[8]),
    .o(al_cbbf04f9));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*B*~A)"),
    .INIT(64'h0000000000000004))
    al_15d7a978 (
    .a(al_8afe6a9f),
    .b(al_cbbf04f9),
    .c(al_821706b3[0]),
    .d(al_821706b3[1]),
    .e(al_821706b3[2]),
    .f(al_821706b3[3]),
    .o(al_1e8f68ca));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(A*(B*D*~(E)+~(B)*~(D)*E)))"),
    .INIT(32'h0f0d070f))
    al_71d17667 (
    .a(al_1e8f68ca),
    .b(al_edc29fee),
    .c(al_e199650d),
    .d(al_821706b3[6]),
    .e(al_821706b3[9]),
    .o(al_75356484));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(~D*B)))"),
    .INIT(16'h0545))
    al_7f79fad (
    .a(al_75356484),
    .b(al_8f22b7e0),
    .c(al_33f2071f),
    .d(al_c925873),
    .o(al_bb3ef93c));
  AL_MAP_LUT6 #(
    .EQN("(~(~D*C)*~(F*E*~(B*A)))"),
    .INIT(64'h8808ff0fff0fff0f))
    al_db1e9dd (
    .a(al_2337d80f),
    .b(al_87969af9),
    .c(al_85bba154),
    .d(al_a494216e),
    .e(al_1d8c2b07),
    .f(al_4fb6999c),
    .o(al_5227328));
  AL_MAP_LUT6 #(
    .EQN("~(A*~(F*E*~(~D*~(C*~B))))"),
    .INIT(64'hff75555555555555))
    al_74db0ee2 (
    .a(al_5227328),
    .b(al_8f22b7e0),
    .c(al_c52cf3e8),
    .d(al_fdd1f60e),
    .e(al_e3f5d0d6),
    .f(al_c35ead5c),
    .o(al_1d84107f));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    al_50d4af44 (
    .a(al_85bba154),
    .b(al_a494216e),
    .c(al_33f2071f),
    .o(al_1491ad5));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    al_e3d5bfa1 (
    .a(al_531ee03c),
    .b(al_33f2071f),
    .c(al_177c7491),
    .d(al_e396ca5d),
    .o(al_aa6ddd9b));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    al_f42e74e7 (
    .a(al_177c7491),
    .b(al_7fe117d0),
    .c(al_5b769262),
    .d(al_72403be8),
    .o(al_4e7d0870));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_d9ecbd21 (
    .a(al_7fe117d0),
    .b(al_5b769262),
    .o(al_964d579));
  AL_MAP_LUT5 #(
    .EQN("(~(~C*~B)*~(E*~(~D*A)))"),
    .INIT(32'h00a8fcfc))
    al_14dfcb43 (
    .a(al_8f22b7e0),
    .b(al_6fa8f988),
    .c(al_c52cf3e8),
    .d(al_ea30f787),
    .e(al_4a548f7c),
    .o(al_32b11a18));
  AL_MAP_LUT6 #(
    .EQN("(~D*~C*~(~B*~A*~(~F*E)))"),
    .INIT(64'h000e000e000f000e))
    al_19382ada (
    .a(al_32b11a18),
    .b(al_20a6f635),
    .c(al_fdd1f60e),
    .d(al_cbafc250),
    .e(al_be1d3817),
    .f(al_4a548f7c),
    .o(al_397de144));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_2be188ef (
    .a(al_e5fcf9b1),
    .b(al_e4dc5a7[0]),
    .o(al_b3c5207a));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_f8e7287f (
    .a(al_eb5c4882),
    .b(al_4d46dbf7[0]),
    .o(al_224d6023[0]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_c99eba5c (
    .a(al_eb5c4882),
    .b(al_4d46dbf7[1]),
    .o(al_224d6023[1]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_8bed3abe (
    .a(al_eb5c4882),
    .b(al_4d46dbf7[2]),
    .o(al_224d6023[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_d713c269 (
    .a(al_eb5c4882),
    .b(al_4d46dbf7[3]),
    .o(al_224d6023[3]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_6de92630 (
    .a(al_eb5c4882),
    .b(al_4d46dbf7[4]),
    .o(al_224d6023[4]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_327f7b3a (
    .a(al_eb5c4882),
    .b(al_4d46dbf7[5]),
    .o(al_224d6023[5]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_477a6285 (
    .a(al_eb5c4882),
    .b(al_4d46dbf7[6]),
    .o(al_224d6023[6]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_348b8dc (
    .a(al_f52ae365),
    .b(al_eb5c4882),
    .c(al_4d46dbf7[7]),
    .o(al_224d6023[7]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C)*~((~B*~A))+D*C*~((~B*~A))+~(D)*C*(~B*~A)+D*C*(~B*~A))"),
    .INIT(16'hfe10))
    al_ed18e1f8 (
    .a(al_b348c1a2),
    .b(al_e2a3cd9),
    .c(al_d75651de),
    .d(al_9affd881[0]),
    .o(al_93cc3d71[0]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C)*~((~B*~A))+D*C*~((~B*~A))+~(D)*C*(~B*~A)+D*C*(~B*~A))"),
    .INIT(16'hfe10))
    al_cea4c138 (
    .a(al_b348c1a2),
    .b(al_e2a3cd9),
    .c(al_d75651de),
    .d(al_9affd881[1]),
    .o(al_93cc3d71[1]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C)*~((~B*~A))+D*C*~((~B*~A))+~(D)*C*(~B*~A)+D*C*(~B*~A))"),
    .INIT(16'hfe10))
    al_a90b8cab (
    .a(al_b348c1a2),
    .b(al_e2a3cd9),
    .c(al_d75651de),
    .d(al_9affd881[2]),
    .o(al_93cc3d71[2]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C)*~((~B*~A))+D*C*~((~B*~A))+~(D)*C*(~B*~A)+D*C*(~B*~A))"),
    .INIT(16'hfe10))
    al_f085f2a7 (
    .a(al_b348c1a2),
    .b(al_e2a3cd9),
    .c(al_d75651de),
    .d(al_9affd881[3]),
    .o(al_93cc3d71[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    al_26194053 (
    .a(al_b348c1a2),
    .b(al_e2a3cd9),
    .c(al_9affd881[4]),
    .o(al_93cc3d71[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    al_7aa2334f (
    .a(al_b348c1a2),
    .b(al_e2a3cd9),
    .c(al_9affd881[5]),
    .o(al_93cc3d71[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    al_aa0795e5 (
    .a(al_b348c1a2),
    .b(al_e2a3cd9),
    .c(al_9affd881[6]),
    .o(al_93cc3d71[6]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    al_ebb56842 (
    .a(al_b348c1a2),
    .b(al_e2a3cd9),
    .c(al_9affd881[7]),
    .o(al_93cc3d71[7]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_8ec76144 (
    .a(al_e5fcf9b1),
    .b(al_84c0beb4[0]),
    .o(al_9595c97a[0]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_af580c11 (
    .a(al_e5fcf9b1),
    .b(al_84c0beb4[1]),
    .o(al_9595c97a[1]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_fc6355b (
    .a(al_e5fcf9b1),
    .b(al_84c0beb4[2]),
    .o(al_9595c97a[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_efade4f5 (
    .a(al_e5fcf9b1),
    .b(al_84c0beb4[3]),
    .o(al_9595c97a[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_75082a4e (
    .a(al_e5fcf9b1),
    .b(al_84c0beb4[4]),
    .o(al_9595c97a[4]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_6a695af8 (
    .a(al_e5fcf9b1),
    .b(al_84c0beb4[5]),
    .o(al_9595c97a[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_d6aaa21c (
    .a(al_e5fcf9b1),
    .b(al_84c0beb4[6]),
    .o(al_9595c97a[6]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_875015c2 (
    .a(al_e5fcf9b1),
    .b(al_84c0beb4[7]),
    .o(al_9595c97a[7]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_cf61a839 (
    .a(al_72403be8),
    .b(al_643ac1f2),
    .c(al_68ba43d4),
    .o(al_d277135));
  AL_MAP_LUT4 #(
    .EQN("~(~C*A*~(D*~B))"),
    .INIT(16'hf7f5))
    al_461148f2 (
    .a(al_8f22b7e0),
    .b(al_c52cf3e8),
    .c(al_cbafc250),
    .d(al_c925873),
    .o(al_f28fd6dc));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*~A)"),
    .INIT(16'h0040))
    al_7fbdae39 (
    .a(al_1698ebe9),
    .b(al_e3f5d0d6),
    .c(al_c35ead5c),
    .d(al_f28e4921),
    .o(al_567fa47e));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(E*~D*~C*B))"),
    .INIT(32'haaaeaaaa))
    al_34f0bb0f (
    .a(al_567fa47e),
    .b(al_d1e17be4),
    .c(al_edc29fee),
    .d(al_177c7491),
    .e(al_f28e4921),
    .o(al_7f7f4148));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(~D*~A))"),
    .INIT(16'h0302))
    al_e9e6a2b4 (
    .a(al_279c902b),
    .b(al_206f470e),
    .c(al_f28e4921),
    .d(al_21d722fe),
    .o(al_ab82ee9a));
  AL_MAP_LUT6 #(
    .EQN("(~E*~D*~(~F*~(A*~(~C*B))))"),
    .INIT(64'h000000ff000000a2))
    al_73b45bb5 (
    .a(al_279c902b),
    .b(al_4ba3ac36),
    .c(al_33f2071f),
    .d(al_206f470e),
    .e(al_f28e4921),
    .f(al_b65fd623),
    .o(al_95d27a4c));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_5cfbaccd (
    .a(al_ee74aec5),
    .b(al_b984f6c1),
    .c(al_bc147132),
    .o(al_2337d80f));
  AL_MAP_LUT6 #(
    .EQN("(D*C*~(B*~(~F*~(~E*A))))"),
    .INIT(64'h30003000f0007000))
    al_eab229f9 (
    .a(al_2e2debcb),
    .b(al_cbafc250),
    .c(al_1d8c2b07),
    .d(al_4fb6999c),
    .e(al_5f257019[5]),
    .f(al_e199650d),
    .o(al_1dbbddf2));
  AL_MAP_LUT6 #(
    .EQN("~(~(~F*E)*~(C*B*~(~D*~A)))"),
    .INIT(64'hc080c080ffffc080))
    al_f510af6b (
    .a(al_1dbbddf2),
    .b(al_2337d80f),
    .c(al_87969af9),
    .d(al_85bba154),
    .e(al_a494216e),
    .f(al_33f2071f),
    .o(al_af806095));
  AL_MAP_LUT4 #(
    .EQN("~(~(~C*B)*~(D*~A))"),
    .INIT(16'h5d0c))
    al_1dc0b5cb (
    .a(al_33f2071f),
    .b(al_13f48428),
    .c(al_b65fd623),
    .d(al_2b1074ba),
    .o(al_8aeddbc));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*A)"),
    .INIT(64'h8000000000000000))
    al_52d9f39f (
    .a(al_1bfb1d64),
    .b(al_af1ac2b6),
    .c(al_75182ad3),
    .d(al_5ad7d7e7),
    .e(al_c5664b3b),
    .f(al_9f6ea2ef),
    .o(al_8f0a5b42));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_e15b003f (
    .a(al_8f0a5b42),
    .b(al_ad4aba0),
    .o(al_cafc0d92));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_13a263c9 (
    .a(al_33f2071f),
    .b(al_177c7491),
    .o(al_db73eae9));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*~B*~(~D*~C)))"),
    .INIT(32'haaaa888a))
    al_20163cd4 (
    .a(al_a494216e),
    .b(al_77192586),
    .c(al_e702d1c[0]),
    .d(al_e702d1c[1]),
    .e(al_e702d1c[2]),
    .o(al_97576f4d));
  AL_MAP_LUT6 #(
    .EQN("~(~A*~(~E*~(~C*~(F*D*B))))"),
    .INIT(64'haaaafefaaaaafafa))
    al_15f33769 (
    .a(al_97576f4d),
    .b(al_8f22b7e0),
    .c(al_db73eae9),
    .d(al_c52cf3e8),
    .e(al_cbafc250),
    .f(al_c35ead5c),
    .o(al_64c768d));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(A)*~(D)+~(~C*~B)*A*~(D)+~(~(~C*~B))*A*D+~(~C*~B)*A*D)"),
    .INIT(16'haafc))
    al_c5282146 (
    .a(al_64fd2ef5[0]),
    .b(al_efc7f78a[0]),
    .c(al_efc7f78a[14]),
    .d(al_25d4a5f3),
    .o(al_ecab3deb[0]));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(A)*~(D)+~(~C*~B)*A*~(D)+~(~(~C*~B))*A*D+~(~C*~B)*A*D)"),
    .INIT(16'haafc))
    al_4a0e1470 (
    .a(al_64fd2ef5[10]),
    .b(al_efc7f78a[10]),
    .c(al_efc7f78a[14]),
    .d(al_25d4a5f3),
    .o(al_ecab3deb[10]));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(A)*~(D)+~(~C*~B)*A*~(D)+~(~(~C*~B))*A*D+~(~C*~B)*A*D)"),
    .INIT(16'haafc))
    al_372757a8 (
    .a(al_64fd2ef5[11]),
    .b(al_efc7f78a[11]),
    .c(al_efc7f78a[14]),
    .d(al_25d4a5f3),
    .o(al_ecab3deb[11]));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(A)*~(D)+~(~C*~B)*A*~(D)+~(~(~C*~B))*A*D+~(~C*~B)*A*D)"),
    .INIT(16'haafc))
    al_427f07cf (
    .a(al_64fd2ef5[12]),
    .b(al_efc7f78a[12]),
    .c(al_efc7f78a[14]),
    .d(al_25d4a5f3),
    .o(al_ecab3deb[12]));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(A)*~(D)+~(~C*~B)*A*~(D)+~(~(~C*~B))*A*D+~(~C*~B)*A*D)"),
    .INIT(16'haafc))
    al_9d450f27 (
    .a(al_64fd2ef5[13]),
    .b(al_efc7f78a[13]),
    .c(al_efc7f78a[14]),
    .d(al_25d4a5f3),
    .o(al_ecab3deb[13]));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(A)*~(D)+~(~C*~B)*A*~(D)+~(~(~C*~B))*A*D+~(~C*~B)*A*D)"),
    .INIT(16'haafc))
    al_5e04eeff (
    .a(al_64fd2ef5[1]),
    .b(al_efc7f78a[1]),
    .c(al_efc7f78a[14]),
    .d(al_25d4a5f3),
    .o(al_ecab3deb[1]));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(A)*~(D)+~(~C*~B)*A*~(D)+~(~(~C*~B))*A*D+~(~C*~B)*A*D)"),
    .INIT(16'haafc))
    al_cfedf04b (
    .a(al_64fd2ef5[2]),
    .b(al_efc7f78a[2]),
    .c(al_efc7f78a[14]),
    .d(al_25d4a5f3),
    .o(al_ecab3deb[2]));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(A)*~(D)+~(~C*~B)*A*~(D)+~(~(~C*~B))*A*D+~(~C*~B)*A*D)"),
    .INIT(16'haafc))
    al_f2d88db (
    .a(al_64fd2ef5[3]),
    .b(al_efc7f78a[3]),
    .c(al_efc7f78a[14]),
    .d(al_25d4a5f3),
    .o(al_ecab3deb[3]));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(A)*~(D)+~(~C*~B)*A*~(D)+~(~(~C*~B))*A*D+~(~C*~B)*A*D)"),
    .INIT(16'haafc))
    al_c19fb52c (
    .a(al_64fd2ef5[4]),
    .b(al_efc7f78a[4]),
    .c(al_efc7f78a[14]),
    .d(al_25d4a5f3),
    .o(al_ecab3deb[4]));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(A)*~(D)+~(~C*~B)*A*~(D)+~(~(~C*~B))*A*D+~(~C*~B)*A*D)"),
    .INIT(16'haafc))
    al_2f6b875f (
    .a(al_64fd2ef5[5]),
    .b(al_efc7f78a[5]),
    .c(al_efc7f78a[14]),
    .d(al_25d4a5f3),
    .o(al_ecab3deb[5]));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(A)*~(D)+~(~C*~B)*A*~(D)+~(~(~C*~B))*A*D+~(~C*~B)*A*D)"),
    .INIT(16'haafc))
    al_9acfbd60 (
    .a(al_64fd2ef5[6]),
    .b(al_efc7f78a[6]),
    .c(al_efc7f78a[14]),
    .d(al_25d4a5f3),
    .o(al_ecab3deb[6]));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(A)*~(D)+~(~C*~B)*A*~(D)+~(~(~C*~B))*A*D+~(~C*~B)*A*D)"),
    .INIT(16'haafc))
    al_bfa7a6a0 (
    .a(al_64fd2ef5[7]),
    .b(al_efc7f78a[7]),
    .c(al_efc7f78a[14]),
    .d(al_25d4a5f3),
    .o(al_ecab3deb[7]));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(A)*~(D)+~(~C*~B)*A*~(D)+~(~(~C*~B))*A*D+~(~C*~B)*A*D)"),
    .INIT(16'haafc))
    al_70beeb38 (
    .a(al_64fd2ef5[8]),
    .b(al_efc7f78a[8]),
    .c(al_efc7f78a[14]),
    .d(al_25d4a5f3),
    .o(al_ecab3deb[8]));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*~B)*~(A)*~(D)+~(~C*~B)*A*~(D)+~(~(~C*~B))*A*D+~(~C*~B)*A*D)"),
    .INIT(16'haafc))
    al_3405b1e0 (
    .a(al_64fd2ef5[9]),
    .b(al_efc7f78a[9]),
    .c(al_efc7f78a[14]),
    .d(al_25d4a5f3),
    .o(al_ecab3deb[9]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*~A))"),
    .INIT(8'hdc))
    al_ee54219e (
    .a(al_33f2071f),
    .b(al_643ac1f2),
    .c(al_25d4a5f3),
    .o(al_8b965f41));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*~D)*~(~C*B*A))"),
    .INIT(32'h08ff0808))
    al_d7d4883a (
    .a(al_2e2debcb),
    .b(al_cbafc250),
    .c(al_5f257019[5]),
    .d(al_f28e4921),
    .e(al_4dac203f),
    .o(al_66382828));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~C)*~(B*~A))"),
    .INIT(16'h4f44))
    al_8eacac3e (
    .a(al_13f48428),
    .b(al_3e886516),
    .c(al_f28e4921),
    .d(al_6980bc30),
    .o(al_5156ba29));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    al_1013c70f (
    .a(al_24ac8493[0]),
    .b(al_24ac8493[1]),
    .c(al_24ac8493[2]),
    .d(al_eb5c4882),
    .o(al_1a33f9b0));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*(~C*B)*~(D)*~(E)+A*(~C*B)*~(D)*~(E)+~(A)*~((~C*B))*~(D)*E+A*~((~C*B))*~(D)*E+~(A)*(~C*B)*~(D)*E+A*(~C*B)*~(D)*E+~(A)*~((~C*B))*D*E)"),
    .INIT(32'h51ff000c))
    al_d01443a3 (
    .a(al_1a33f9b0),
    .b(al_2337d80f),
    .c(al_9a8c459a),
    .d(al_f92026f1),
    .e(al_a978a29f),
    .o(al_4854aa2f));
  AL_MAP_LUT5 #(
    .EQN("(~(~D*~C)*~(E*~B*A))"),
    .INIT(32'hddd0fff0))
    al_66c3c13c (
    .a(al_33f2071f),
    .b(al_c925873),
    .c(al_f28e4921),
    .d(al_3475fb1c),
    .e(al_beea368e),
    .o(al_5cd49131));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    al_224097bc (
    .a(al_8aa33695),
    .b(al_5cd49131),
    .c(al_a978a29f),
    .o(al_e03ae0c1));
  AL_MAP_LUT4 #(
    .EQN("(A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'ha280))
    al_cf8b8215 (
    .a(al_d1e17be4),
    .b(al_177c7491),
    .c(al_3475fb1c),
    .d(al_8b86ece7),
    .o(al_508b6c4c));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_f2e43996 (
    .a(al_d1e17be4),
    .b(al_a494216e),
    .c(al_e20fd0c7[0]),
    .o(al_4b4b7bbc[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_c2333c62 (
    .a(al_d1e17be4),
    .b(al_a494216e),
    .c(al_e20fd0c7[10]),
    .o(al_4b4b7bbc[10]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*A)"),
    .INIT(8'hf7))
    al_79d8ceac (
    .a(al_d1e17be4),
    .b(al_a494216e),
    .c(al_e20fd0c7[11]),
    .o(al_4b4b7bbc[11]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_7c5b99ad (
    .a(al_d1e17be4),
    .b(al_a494216e),
    .c(al_e20fd0c7[12]),
    .o(al_4b4b7bbc[12]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_6061b9bc (
    .a(al_d1e17be4),
    .b(al_a494216e),
    .c(al_e20fd0c7[13]),
    .o(al_4b4b7bbc[13]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D)*~((C*A))+~B*D*~((C*A))+~(~B)*D*(C*A)+~B*D*(C*A))"),
    .INIT(16'hb313))
    al_5ef58975 (
    .a(al_d1e17be4),
    .b(al_edc29fee),
    .c(al_a494216e),
    .d(al_e20fd0c7[14]),
    .o(al_4b4b7bbc[14]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_27c3d7e4 (
    .a(al_d1e17be4),
    .b(al_a494216e),
    .c(al_e20fd0c7[1]),
    .o(al_4b4b7bbc[1]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*A)"),
    .INIT(8'hf7))
    al_a118d03f (
    .a(al_d1e17be4),
    .b(al_a494216e),
    .c(al_e20fd0c7[2]),
    .o(al_4b4b7bbc[2]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D)*~((C*A))+~B*D*~((C*A))+~(~B)*D*(C*A)+~B*D*(C*A))"),
    .INIT(16'hb313))
    al_6cfedb7d (
    .a(al_d1e17be4),
    .b(al_edc29fee),
    .c(al_a494216e),
    .d(al_e20fd0c7[3]),
    .o(al_4b4b7bbc[3]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D)*~((C*A))+B*D*~((C*A))+~(B)*D*(C*A)+B*D*(C*A))"),
    .INIT(16'hec4c))
    al_6ccafe52 (
    .a(al_d1e17be4),
    .b(al_edc29fee),
    .c(al_a494216e),
    .d(al_e20fd0c7[4]),
    .o(al_4b4b7bbc[4]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D)*~((C*A))+~B*D*~((C*A))+~(~B)*D*(C*A)+~B*D*(C*A))"),
    .INIT(16'hb313))
    al_76dad919 (
    .a(al_d1e17be4),
    .b(al_edc29fee),
    .c(al_a494216e),
    .d(al_e20fd0c7[5]),
    .o(al_4b4b7bbc[5]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*A)"),
    .INIT(8'hf7))
    al_6aaead76 (
    .a(al_d1e17be4),
    .b(al_a494216e),
    .c(al_e20fd0c7[6]),
    .o(al_4b4b7bbc[6]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*A)"),
    .INIT(8'hf7))
    al_fa24b654 (
    .a(al_d1e17be4),
    .b(al_a494216e),
    .c(al_e20fd0c7[7]),
    .o(al_4b4b7bbc[7]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*A)"),
    .INIT(8'hf7))
    al_5bca2c77 (
    .a(al_d1e17be4),
    .b(al_a494216e),
    .c(al_e20fd0c7[8]),
    .o(al_4b4b7bbc[8]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*A)"),
    .INIT(8'hf7))
    al_626a3459 (
    .a(al_d1e17be4),
    .b(al_a494216e),
    .c(al_e20fd0c7[9]),
    .o(al_4b4b7bbc[9]));
  AL_MAP_LUT6 #(
    .EQN("~(~(~F*E*~C*B)*~(D*A))"),
    .INIT(64'haa00aa00ae0caa00))
    al_80272635 (
    .a(al_e1420a1f),
    .b(al_531ee03c),
    .c(al_a494216e),
    .d(al_33f2071f),
    .e(al_177c7491),
    .f(al_cbafc250),
    .o(al_acdc1781));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_8495cfe0 (
    .a(al_8e462c61[0]),
    .b(al_8e462c61[1]),
    .c(al_8e462c61[2]),
    .d(al_8e462c61[3]),
    .o(al_1638f286));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    al_6320cb28 (
    .a(al_1638f286),
    .b(al_8e462c61[4]),
    .c(al_8e462c61[5]),
    .d(al_8e462c61[6]),
    .e(al_8e462c61[7]),
    .o(al_44b2d585));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_38e94faa (
    .a(al_8e462c61[8]),
    .b(al_8e462c61[9]),
    .c(al_8e462c61[10]),
    .d(al_8e462c61[11]),
    .o(al_6b4822fe));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    al_bdbc8f3 (
    .a(al_44b2d585),
    .b(al_6b4822fe),
    .c(al_8e462c61[12]),
    .d(al_8e462c61[13]),
    .e(al_8e462c61[14]),
    .o(al_fc7de59c));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*~B))"),
    .INIT(8'hba))
    al_bd965852 (
    .a(al_fc7de59c),
    .b(al_f28e4921),
    .c(al_d224660a),
    .o(al_4d4a65fe));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_a5e64ccf (
    .a(al_ecd47e95),
    .b(al_821706b3[0]),
    .o(al_93f1315e[0]));
  AL_MAP_LUT3 #(
    .EQN("(~A*(C@B))"),
    .INIT(8'h14))
    al_60e1e274 (
    .a(al_ecd47e95),
    .b(al_821706b3[0]),
    .c(al_821706b3[1]),
    .o(al_93f1315e[1]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D@(C*B)))"),
    .INIT(16'h1540))
    al_86e5dc4c (
    .a(al_ecd47e95),
    .b(al_821706b3[0]),
    .c(al_821706b3[1]),
    .d(al_821706b3[2]),
    .o(al_93f1315e[2]));
  AL_MAP_LUT5 #(
    .EQN("(~A*(E@(D*C*B)))"),
    .INIT(32'h15554000))
    al_d442a8a4 (
    .a(al_ecd47e95),
    .b(al_821706b3[0]),
    .c(al_821706b3[1]),
    .d(al_821706b3[2]),
    .e(al_821706b3[3]),
    .o(al_93f1315e[3]));
  AL_MAP_LUT6 #(
    .EQN("(~A*(F@(E*D*C*B)))"),
    .INIT(64'h1555555540000000))
    al_95746355 (
    .a(al_ecd47e95),
    .b(al_821706b3[0]),
    .c(al_821706b3[1]),
    .d(al_821706b3[2]),
    .e(al_821706b3[3]),
    .f(al_821706b3[4]),
    .o(al_93f1315e[4]));
  AL_MAP_LUT6 #(
    .EQN("(F@(E*D*C*B*A))"),
    .INIT(64'h7fffffff80000000))
    al_18b19a9c (
    .a(al_821706b3[0]),
    .b(al_821706b3[1]),
    .c(al_821706b3[2]),
    .d(al_821706b3[3]),
    .e(al_821706b3[4]),
    .f(al_821706b3[5]),
    .o(al_dcce7f97[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_f884e27e (
    .a(al_ecd47e95),
    .b(al_dcce7f97[5]),
    .o(al_93f1315e[5]));
  AL_MAP_LUT3 #(
    .EQN("(~A*(C@B))"),
    .INIT(8'h14))
    al_14f4de4a (
    .a(al_ecd47e95),
    .b(al_f51408c3),
    .c(al_821706b3[6]),
    .o(al_93f1315e[6]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D@(C*B)))"),
    .INIT(16'h1540))
    al_452253fb (
    .a(al_ecd47e95),
    .b(al_f51408c3),
    .c(al_821706b3[6]),
    .d(al_821706b3[7]),
    .o(al_93f1315e[7]));
  AL_MAP_LUT5 #(
    .EQN("(~A*(E@(D*C*B)))"),
    .INIT(32'h15554000))
    al_1da2eda (
    .a(al_ecd47e95),
    .b(al_f51408c3),
    .c(al_821706b3[6]),
    .d(al_821706b3[7]),
    .e(al_821706b3[8]),
    .o(al_93f1315e[8]));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*A)"),
    .INIT(64'h8000000000000000))
    al_3f651589 (
    .a(al_821706b3[0]),
    .b(al_821706b3[1]),
    .c(al_821706b3[2]),
    .d(al_821706b3[3]),
    .e(al_821706b3[4]),
    .f(al_821706b3[5]),
    .o(al_f51408c3));
  AL_MAP_LUT6 #(
    .EQN("(~A*(F@(E*D*C*B)))"),
    .INIT(64'h1555555540000000))
    al_4ef4ebc4 (
    .a(al_ecd47e95),
    .b(al_f51408c3),
    .c(al_821706b3[6]),
    .d(al_821706b3[7]),
    .e(al_821706b3[8]),
    .f(al_821706b3[9]),
    .o(al_93f1315e[9]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D@(~B*~A)))"),
    .INIT(16'h10e0))
    al_6d23823f (
    .a(al_1f250659),
    .b(al_8aa33695),
    .c(al_1104f08c),
    .d(al_8c490204[0]),
    .o(al_c8474427[0]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_8c0649ea (
    .a(al_8c490204[0]),
    .b(al_8c490204[1]),
    .c(al_8c490204[2]),
    .d(al_8c490204[3]),
    .o(al_c91a5908));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    al_b84d175 (
    .a(al_c91a5908),
    .b(al_8c490204[4]),
    .c(al_8c490204[5]),
    .d(al_8c490204[6]),
    .e(al_8c490204[7]),
    .o(al_7fb47a00));
  AL_MAP_LUT5 #(
    .EQN("(E*A*~(D*~C*~B))"),
    .INIT(32'ha8aa0000))
    al_777abe9a (
    .a(al_7fb47a00),
    .b(al_b156040b),
    .c(al_8aa33695),
    .d(al_51172105),
    .e(al_8c490204[8]),
    .o(al_900fca1b));
  AL_MAP_LUT4 #(
    .EQN("(B*(D@(C*A)))"),
    .INIT(16'h4c80))
    al_cd3b039e (
    .a(al_900fca1b),
    .b(al_1104f08c),
    .c(al_8c490204[9]),
    .d(al_8c490204[10]),
    .o(al_c8474427[10]));
  AL_MAP_LUT5 #(
    .EQN("(C*(E@(D*~(~B*~A))))"),
    .INIT(32'h10f0e000))
    al_75cabd28 (
    .a(al_1f250659),
    .b(al_8aa33695),
    .c(al_1104f08c),
    .d(al_8c490204[0]),
    .e(al_8c490204[1]),
    .o(al_c8474427[1]));
  AL_MAP_LUT6 #(
    .EQN("(C*(F@(E*D*~(~B*~A))))"),
    .INIT(64'h10f0f0f0e0000000))
    al_a5216ff0 (
    .a(al_1f250659),
    .b(al_8aa33695),
    .c(al_1104f08c),
    .d(al_8c490204[0]),
    .e(al_8c490204[1]),
    .f(al_8c490204[2]),
    .o(al_c8474427[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_909162b0 (
    .a(al_8c490204[0]),
    .b(al_8c490204[1]),
    .c(al_8c490204[2]),
    .o(al_5b8b9ce6));
  AL_MAP_LUT5 #(
    .EQN("(C*(E@(D*~(~B*~A))))"),
    .INIT(32'h10f0e000))
    al_5470c403 (
    .a(al_1f250659),
    .b(al_8aa33695),
    .c(al_1104f08c),
    .d(al_5b8b9ce6),
    .e(al_8c490204[3]),
    .o(al_c8474427[3]));
  AL_MAP_LUT3 #(
    .EQN("(B*(C@A))"),
    .INIT(8'h48))
    al_3566c3b8 (
    .a(al_d9ca5f64),
    .b(al_1104f08c),
    .c(al_8c490204[4]),
    .o(al_c8474427[4]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D@(C*A)))"),
    .INIT(16'h4c80))
    al_edf7a082 (
    .a(al_d9ca5f64),
    .b(al_1104f08c),
    .c(al_8c490204[4]),
    .d(al_8c490204[5]),
    .o(al_c8474427[5]));
  AL_MAP_LUT5 #(
    .EQN("(B*(E@(D*C*A)))"),
    .INIT(32'h4ccc8000))
    al_8e2f0c75 (
    .a(al_d9ca5f64),
    .b(al_1104f08c),
    .c(al_8c490204[4]),
    .d(al_8c490204[5]),
    .e(al_8c490204[6]),
    .o(al_c8474427[6]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*~A))"),
    .INIT(16'hef00))
    al_c942164e (
    .a(al_b156040b),
    .b(al_8aa33695),
    .c(al_51172105),
    .d(al_c91a5908),
    .o(al_d9ca5f64));
  AL_MAP_LUT6 #(
    .EQN("(B*(F@(E*D*C*A)))"),
    .INIT(64'h4ccccccc80000000))
    al_a14937b1 (
    .a(al_d9ca5f64),
    .b(al_1104f08c),
    .c(al_8c490204[4]),
    .d(al_8c490204[5]),
    .e(al_8c490204[6]),
    .f(al_8c490204[7]),
    .o(al_c8474427[7]));
  AL_MAP_LUT5 #(
    .EQN("(D*(E@(B*~(~C*~A))))"),
    .INIT(32'h3700c800))
    al_e52fce44 (
    .a(al_1f250659),
    .b(al_7fb47a00),
    .c(al_8aa33695),
    .d(al_1104f08c),
    .e(al_8c490204[8]),
    .o(al_c8474427[8]));
  AL_MAP_LUT3 #(
    .EQN("(B*(C@A))"),
    .INIT(8'h48))
    al_aa7e8612 (
    .a(al_900fca1b),
    .b(al_1104f08c),
    .c(al_8c490204[9]),
    .o(al_c8474427[9]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    al_823c1e1f (
    .a(al_d1e17be4),
    .b(al_edc29fee),
    .c(al_85bba154),
    .d(al_a494216e),
    .e(al_cbafc250),
    .o(al_1104f08c));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_6e386b0c (
    .a(al_8c490204[5]),
    .b(al_8c490204[6]),
    .c(al_8c490204[7]),
    .d(al_8c490204[8]),
    .o(al_3cdb7f2c));
  AL_MAP_LUT6 #(
    .EQN("(F*~(~E*~D*A*~(C*B)))"),
    .INIT(64'hffffffd500000000))
    al_ca6ff5cd (
    .a(al_3cdb7f2c),
    .b(al_8c490204[1]),
    .c(al_8c490204[2]),
    .d(al_8c490204[3]),
    .e(al_8c490204[4]),
    .f(al_8c490204[9]),
    .o(al_ee9e22e));
  AL_MAP_LUT5 #(
    .EQN("(~(D*~C*~B)*~(~E*~A))"),
    .INIT(32'hfcffa8aa))
    al_86526535 (
    .a(al_ee9e22e),
    .b(al_b156040b),
    .c(al_8aa33695),
    .d(al_51172105),
    .e(al_8c490204[10]),
    .o(al_addc1415));
  AL_MAP_LUT5 #(
    .EQN("~(~D*C*~(B*~(~E*~A)))"),
    .INIT(32'hffcfff8f))
    al_365121a (
    .a(al_addc1415),
    .b(al_1104f08c),
    .c(al_d1e17be4),
    .d(al_edc29fee),
    .e(al_4a548f7c),
    .o(al_f2d6f40b));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E*~D*~C*~B))"),
    .INIT(32'h55545555))
    al_75ae302c (
    .a(al_33f2071f),
    .b(al_cbafc250),
    .c(al_1d8c2b07),
    .d(al_b7729dd8),
    .e(al_77192586),
    .o(al_756a1d77));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_b9134511 (
    .a(al_756a1d77),
    .b(al_d1e17be4),
    .c(al_edc29fee),
    .o(al_81aa4d04));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    al_9a6f60f0 (
    .a(al_7fe117d0),
    .b(al_5b769262),
    .c(al_72403be8),
    .d(al_cbafc250),
    .o(al_d6cf9565));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(~E*D*~(~C*B)))"),
    .INIT(32'haaaafbaa))
    al_a65c79 (
    .a(al_d6cf9565),
    .b(al_2337d80f),
    .c(al_279c902b),
    .d(al_177c7491),
    .e(al_643ac1f2),
    .o(al_ab89cd63));
  AL_DFF_X al_d509de0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_ifg_val[0]),
    .en(al_520be21e),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_984d3b84[0]));
  AL_DFF_X al_6ddac1c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_ifg_val[1]),
    .en(al_520be21e),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_984d3b84[1]));
  AL_DFF_X al_6a5fbea5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_ifg_val[2]),
    .en(al_520be21e),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_984d3b84[2]));
  AL_DFF_X al_f637b416 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_ifg_val[3]),
    .en(al_520be21e),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_984d3b84[3]));
  AL_DFF_X al_55487ece (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_ifg_val[4]),
    .en(al_520be21e),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_984d3b84[4]));
  AL_DFF_X al_80d9aa3e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_ifg_val[5]),
    .en(al_520be21e),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_984d3b84[5]));
  AL_DFF_X al_6ae4c6c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_ifg_val[6]),
    .en(al_520be21e),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_984d3b84[6]));
  AL_DFF_X al_9b24ba4b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(tx_ifg_val[7]),
    .en(al_520be21e),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_984d3b84[7]));
  AL_DFF_X al_b526117d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ae339d26[2]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_19bf88c2[2]));
  AL_DFF_X al_eb81c3da (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d09ba8fa),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_19bf88c2[4]));
  AL_DFF_X al_575064ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5db4ba74[0]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_4d46dbf7[0]));
  AL_DFF_X al_3bfd73dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5db4ba74[1]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_4d46dbf7[1]));
  AL_DFF_X al_d8e6799b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5db4ba74[2]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_4d46dbf7[2]));
  AL_DFF_X al_140a8b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5db4ba74[3]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_4d46dbf7[3]));
  AL_DFF_X al_f8c18f8f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5db4ba74[4]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_4d46dbf7[4]));
  AL_DFF_X al_8e36fb89 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5db4ba74[5]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_4d46dbf7[5]));
  AL_DFF_X al_dcb33971 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5db4ba74[6]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_4d46dbf7[6]));
  AL_DFF_X al_46ad8924 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_5db4ba74[7]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_4d46dbf7[7]));
  AL_DFF_X al_75a2ae36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_224d6023[0]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9affd881[0]));
  AL_DFF_X al_c4e22be8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_224d6023[1]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9affd881[1]));
  AL_DFF_X al_da8e0c62 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_224d6023[2]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9affd881[2]));
  AL_DFF_X al_288224e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_224d6023[3]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9affd881[3]));
  AL_DFF_X al_497cf6e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_224d6023[4]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9affd881[4]));
  AL_DFF_X al_f9a1e727 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_224d6023[5]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9affd881[5]));
  AL_DFF_X al_6dcf5b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_224d6023[6]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9affd881[6]));
  AL_DFF_X al_310e6b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_224d6023[7]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_9affd881[7]));
  AL_DFF_X al_28587a24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_93cc3d71[0]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_84c0beb4[0]));
  AL_DFF_X al_78e87bae (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_93cc3d71[1]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_84c0beb4[1]));
  AL_DFF_X al_a1095b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_93cc3d71[2]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_84c0beb4[2]));
  AL_DFF_X al_dbb18bdb (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_93cc3d71[3]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_84c0beb4[3]));
  AL_DFF_X al_9151909c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_93cc3d71[4]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_84c0beb4[4]));
  AL_DFF_X al_2d603ea8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_93cc3d71[5]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_84c0beb4[5]));
  AL_DFF_X al_14bf1f49 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_93cc3d71[6]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_84c0beb4[6]));
  AL_DFF_X al_495e4b64 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_93cc3d71[7]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_84c0beb4[7]));
  AL_DFF_X al_6415bfdc (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9595c97a[0]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_8a6ca59e[0]));
  AL_DFF_X al_34fe6897 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9595c97a[1]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_8a6ca59e[1]));
  AL_DFF_X al_fd866596 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9595c97a[2]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_8a6ca59e[2]));
  AL_DFF_X al_25b737de (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9595c97a[3]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_8a6ca59e[3]));
  AL_DFF_X al_90281169 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9595c97a[4]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_8a6ca59e[4]));
  AL_DFF_X al_e66208e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9595c97a[5]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_8a6ca59e[5]));
  AL_DFF_X al_ff226a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9595c97a[6]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_8a6ca59e[6]));
  AL_DFF_X al_5a61c6b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9595c97a[7]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_8a6ca59e[7]));
  AL_DFF_X al_8dc26ab6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f83013e9[0]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_e00c8785[0]));
  AL_DFF_X al_b58bcdab (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f83013e9[1]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_e00c8785[1]));
  AL_DFF_X al_40d524af (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f83013e9[2]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_e00c8785[2]));
  AL_DFF_X al_3e7d2466 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f83013e9[3]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_e00c8785[3]));
  AL_DFF_X al_3189625a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f83013e9[4]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_e00c8785[4]));
  AL_DFF_X al_fc5eda39 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f83013e9[5]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_e00c8785[5]));
  AL_DFF_X al_8b452290 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f83013e9[6]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_e00c8785[6]));
  AL_DFF_X al_fa1ab113 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_f83013e9[7]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_e00c8785[7]));
  AL_DFF_X al_a4e4ee24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_48fcd383[8]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_48fcd383[9]));
  AL_DFF_X al_18f09f22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_48fcd383[9]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_48fcd383[10]));
  AL_DFF_X al_fcba3f8a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_48fcd383[10]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_48fcd383[11]));
  AL_DFF_X al_8ccff14c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_48fcd383[11]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_48fcd383[12]));
  AL_DFF_X al_40141f22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_48fcd383[12]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_48fcd383[13]));
  AL_DFF_X al_da2bbb84 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b348c1a2),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_48fcd383[1]));
  AL_DFF_X al_3d967daf (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_48fcd383[1]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_48fcd383[2]));
  AL_DFF_X al_a1ceefea (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_48fcd383[2]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_48fcd383[3]));
  AL_DFF_X al_10181c80 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_48fcd383[3]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_48fcd383[4]));
  AL_DFF_X al_43745815 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_48fcd383[4]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_48fcd383[5]));
  AL_DFF_X al_1486372d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_48fcd383[5]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_48fcd383[6]));
  AL_DFF_X al_2b477cd2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_48fcd383[6]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_48fcd383[7]));
  AL_DFF_X al_8673c959 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_48fcd383[7]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_48fcd383[8]));
  AL_DFF_X al_83511fc4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e2a3cd9),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_e4dc5a7[0]));
  AL_DFF_X al_adbbd817 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e4dc5a7[0]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_e4dc5a7[1]));
  AL_DFF_X al_7f45024f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9affd881[0]),
    .en(al_40a7c639),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_bff87853[0]));
  AL_DFF_X al_8ba5d29d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4d46dbf7[1]),
    .en(al_40a7c639),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_bff87853[9]));
  AL_DFF_X al_afbaf412 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4d46dbf7[2]),
    .en(al_40a7c639),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_bff87853[10]));
  AL_DFF_X al_46fefaf5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4d46dbf7[3]),
    .en(al_40a7c639),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_bff87853[11]));
  AL_DFF_X al_ef384259 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4d46dbf7[4]),
    .en(al_40a7c639),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_bff87853[12]));
  AL_DFF_X al_9306903c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4d46dbf7[5]),
    .en(al_40a7c639),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_bff87853[13]));
  AL_DFF_X al_46f344bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4d46dbf7[6]),
    .en(al_40a7c639),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_bff87853[14]));
  AL_DFF_X al_24f6347f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4d46dbf7[7]),
    .en(al_40a7c639),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_bff87853[15]));
  AL_DFF_X al_4148325d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9affd881[1]),
    .en(al_40a7c639),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_bff87853[1]));
  AL_DFF_X al_80218e37 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9affd881[2]),
    .en(al_40a7c639),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_bff87853[2]));
  AL_DFF_X al_f49cbe46 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9affd881[3]),
    .en(al_40a7c639),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_bff87853[3]));
  AL_DFF_X al_44c5a1af (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9affd881[4]),
    .en(al_40a7c639),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_bff87853[4]));
  AL_DFF_X al_e0ac01a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9affd881[5]),
    .en(al_40a7c639),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_bff87853[5]));
  AL_DFF_X al_48327d5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9affd881[6]),
    .en(al_40a7c639),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_bff87853[6]));
  AL_DFF_X al_821f228e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_9affd881[7]),
    .en(al_40a7c639),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_bff87853[7]));
  AL_DFF_X al_3d5ef7b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4d46dbf7[0]),
    .en(al_40a7c639),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_bff87853[8]));
  AL_DFF_X al_efcfbb60 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_64fd2ef5[0]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_183e87f4[0]));
  AL_DFF_X al_fce0d869 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_64fd2ef5[9]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_183e87f4[9]));
  AL_DFF_X al_7fad46d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_64fd2ef5[10]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_183e87f4[10]));
  AL_DFF_X al_51e790aa (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_64fd2ef5[11]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_183e87f4[11]));
  AL_DFF_X al_bb2e7068 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_64fd2ef5[12]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_183e87f4[12]));
  AL_DFF_X al_888f85dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_64fd2ef5[13]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_183e87f4[13]));
  AL_DFF_X al_152f57b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ecab3deb[0]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_64fd2ef5[0]));
  AL_DFF_X al_1c30fdd6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ecab3deb[1]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_64fd2ef5[1]));
  AL_DFF_X al_63ab1311 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ecab3deb[2]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_64fd2ef5[2]));
  AL_DFF_X al_3ae15d65 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ecab3deb[3]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_64fd2ef5[3]));
  AL_DFF_X al_d050a2ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_64fd2ef5[1]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_183e87f4[1]));
  AL_DFF_X al_f8fdc45 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ecab3deb[4]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_64fd2ef5[4]));
  AL_DFF_X al_cecbfe9a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ecab3deb[5]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_64fd2ef5[5]));
  AL_DFF_X al_b3eba179 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ecab3deb[6]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_64fd2ef5[6]));
  AL_DFF_X al_3e625470 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ecab3deb[7]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_64fd2ef5[7]));
  AL_DFF_X al_3484a07a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ecab3deb[8]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_64fd2ef5[8]));
  AL_DFF_X al_8f63f971 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ecab3deb[9]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_64fd2ef5[9]));
  AL_DFF_X al_be689cfd (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ecab3deb[10]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_64fd2ef5[10]));
  AL_DFF_X al_a19ce700 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ecab3deb[11]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_64fd2ef5[11]));
  AL_DFF_X al_288824d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ecab3deb[12]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_64fd2ef5[12]));
  AL_DFF_X al_59383538 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_ecab3deb[13]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_64fd2ef5[13]));
  AL_DFF_X al_bfc85966 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_64fd2ef5[2]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_183e87f4[2]));
  AL_DFF_X al_b7844ab1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e512aff[0]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_efc7f78a[0]));
  AL_DFF_X al_cc99a2ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e512aff[1]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_efc7f78a[1]));
  AL_DFF_X al_352a2d7f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e512aff[2]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_efc7f78a[2]));
  AL_DFF_X al_1eb849f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e512aff[3]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_efc7f78a[3]));
  AL_DFF_X al_be5f4d39 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e512aff[4]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_efc7f78a[4]));
  AL_DFF_X al_c81335c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e512aff[5]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_efc7f78a[5]));
  AL_DFF_X al_295577bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e512aff[6]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_efc7f78a[6]));
  AL_DFF_X al_9c2d7fcd (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e512aff[7]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_efc7f78a[7]));
  AL_DFF_X al_cbc3de23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e512aff[8]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_efc7f78a[8]));
  AL_DFF_X al_9b1979c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_64fd2ef5[3]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_183e87f4[3]));
  AL_DFF_X al_1bc26213 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e512aff[9]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_efc7f78a[9]));
  AL_DFF_X al_fddc33b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e512aff[10]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_efc7f78a[10]));
  AL_DFF_X al_ed371251 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e512aff[11]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_efc7f78a[11]));
  AL_DFF_X al_c45005f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e512aff[12]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_efc7f78a[12]));
  AL_DFF_X al_ad741cfe (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e512aff[13]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_efc7f78a[13]));
  AL_DFF_X al_deb913f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e512aff[14]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_efc7f78a[14]));
  AL_DFF_X al_3a0de9e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_64fd2ef5[4]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_183e87f4[4]));
  AL_DFF_X al_fdf8b7ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_64fd2ef5[5]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_183e87f4[5]));
  AL_DFF_X al_6d30d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_64fd2ef5[6]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_183e87f4[6]));
  AL_DFF_X al_905493ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_64fd2ef5[7]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_183e87f4[7]));
  AL_DFF_X al_d4495474 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_64fd2ef5[8]),
    .en(al_fbfd813b),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_183e87f4[8]));
  AL_DFF_X al_640f467a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_84a48183[0]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_67d6ec64[0]));
  AL_DFF_X al_851b8c35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_84a48183[1]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_67d6ec64[1]));
  AL_DFF_X al_c2641827 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_84a48183[2]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_67d6ec64[2]));
  AL_DFF_X al_b8d64715 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_84a48183[3]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_67d6ec64[3]));
  AL_DFF_X al_46ecd92c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_84a48183[4]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_67d6ec64[4]));
  AL_DFF_X al_df9cdf27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_84a48183[5]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_67d6ec64[5]));
  AL_DFF_X al_450f7b65 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_84a48183[6]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_67d6ec64[6]));
  AL_DFF_X al_9fc7cf4a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_84a48183[7]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_67d6ec64[7]));
  AL_DFF_X al_f9268aaf (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e23c1f65[0]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_bef8ea23[0]));
  AL_DFF_X al_e48c3d6a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e23c1f65[1]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_bef8ea23[1]));
  AL_DFF_X al_49efc43e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e23c1f65[2]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_bef8ea23[2]));
  AL_DFF_X al_ed76e4fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_e23c1f65[3]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_bef8ea23[3]));
  AL_DFF_X al_903c8b38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4b4b7bbc[0]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_8e462c61[0]));
  AL_DFF_X al_2a2811ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4b4b7bbc[9]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_8e462c61[9]));
  AL_DFF_X al_80da8095 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4b4b7bbc[10]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_8e462c61[10]));
  AL_DFF_X al_8bbc6cdb (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4b4b7bbc[11]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_8e462c61[11]));
  AL_DFF_X al_af0c0e03 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4b4b7bbc[12]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_8e462c61[12]));
  AL_DFF_X al_bb20c936 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4b4b7bbc[13]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_8e462c61[13]));
  AL_DFF_X al_b023207c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4b4b7bbc[14]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_8e462c61[14]));
  AL_DFF_X al_5850995b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4b4b7bbc[1]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_8e462c61[1]));
  AL_DFF_X al_44167216 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4b4b7bbc[2]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_8e462c61[2]));
  AL_DFF_X al_5d479b6f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4b4b7bbc[3]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_8e462c61[3]));
  AL_DFF_X al_65cda8dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4b4b7bbc[4]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_8e462c61[4]));
  AL_DFF_X al_8ca6101f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4b4b7bbc[5]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_8e462c61[5]));
  AL_DFF_X al_b73bbfec (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4b4b7bbc[6]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_8e462c61[6]));
  AL_DFF_X al_afa473a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4b4b7bbc[7]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_8e462c61[7]));
  AL_DFF_X al_81f5fce6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4b4b7bbc[8]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_8e462c61[8]));
  AL_DFF_X al_78016f23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_2b1074ba),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(tx_status_vector[0]));
  AL_DFF_X al_15be4452 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_24da7d44[4]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(tx_status_vector[8]));
  AL_DFF_X al_c55d625f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_24da7d44[5]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(tx_status_vector[9]));
  AL_DFF_X al_f22da1e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_24da7d44[6]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(tx_status_vector[10]));
  AL_DFF_X al_fb14eec7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_24da7d44[7]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(tx_status_vector[11]));
  AL_DFF_X al_386f554a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_24da7d44[8]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(tx_status_vector[12]));
  AL_DFF_X al_f93c11d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_24da7d44[9]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(tx_status_vector[13]));
  AL_DFF_X al_1aa42204 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_24da7d44[10]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(tx_status_vector[14]));
  AL_DFF_X al_1fbea56e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_24da7d44[11]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(tx_status_vector[15]));
  AL_DFF_X al_47182e73 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_24da7d44[12]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(tx_status_vector[16]));
  AL_DFF_X al_c93caeb8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_24da7d44[13]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(tx_status_vector[17]));
  AL_DFF_X al_d1b62ef1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_8f0a5b42),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(tx_status_vector[1]));
  AL_DFF_X al_407a3643 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_19bf88c2[4]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(tx_status_vector[19]));
  AL_DFF_X al_a38acda4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_8b86ece7),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(tx_status_vector[21]));
  AL_DFF_X al_621276f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_d224660a),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(tx_status_vector[22]));
  AL_DFF_X al_5156b6d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_6980bc30),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(tx_status_vector[23]));
  AL_DFF_X al_5ff20413 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4dac203f),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(tx_status_vector[28]));
  AL_DFF_X al_8067bdfe (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_bef8ea23[0]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(tx_status_vector[24]));
  AL_DFF_X al_8bf1b222 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_bef8ea23[1]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(tx_status_vector[25]));
  AL_DFF_X al_5af5a953 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_bef8ea23[2]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(tx_status_vector[26]));
  AL_DFF_X al_6c39f470 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_bef8ea23[3]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(tx_status_vector[27]));
  AL_DFF_X al_65c0e02c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_cafc0d92),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(tx_status_vector[2]));
  AL_DFF_X al_dcad4164 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b65fd623),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(tx_status_vector[20]));
  AL_DFF_X al_d4520540 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_4b2213d6),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(tx_status_vector[18]));
  AL_DFF_X al_debd09fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_24da7d44[0]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(tx_status_vector[4]));
  AL_DFF_X al_d84fdf83 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_24da7d44[1]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(tx_status_vector[5]));
  AL_DFF_X al_4032b87e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_24da7d44[2]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(tx_status_vector[6]));
  AL_DFF_X al_d2cb76d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_24da7d44[3]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(tx_status_vector[7]));
  AL_DFF_X al_5fe64dd0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_93f1315e[0]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_821706b3[0]));
  AL_DFF_X al_5bfe08db (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_93f1315e[9]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_821706b3[9]));
  AL_DFF_X al_1a1e6176 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_93f1315e[1]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_821706b3[1]));
  AL_DFF_X al_e0338f92 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_93f1315e[2]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_821706b3[2]));
  AL_DFF_X al_1fc77a49 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_93f1315e[3]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_821706b3[3]));
  AL_DFF_X al_66c3f19d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_93f1315e[4]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_821706b3[4]));
  AL_DFF_X al_a8bbccef (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_93f1315e[5]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_821706b3[5]));
  AL_DFF_X al_2f0d49cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_93f1315e[6]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_821706b3[6]));
  AL_DFF_X al_6f936a31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_93f1315e[7]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_821706b3[7]));
  AL_DFF_X al_516ca590 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_93f1315e[8]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_821706b3[8]));
  AL_DFF_X al_a7d784b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c8474427[0]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_8c490204[0]));
  AL_DFF_X al_e9596b4c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c8474427[9]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_8c490204[9]));
  AL_DFF_X al_59b21843 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c8474427[10]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_8c490204[10]));
  AL_DFF_X al_1c968819 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c8474427[1]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_8c490204[1]));
  AL_DFF_X al_d6135a30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c8474427[2]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_8c490204[2]));
  AL_DFF_X al_87f934c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c8474427[3]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_8c490204[3]));
  AL_DFF_X al_6bdafb61 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c8474427[4]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_8c490204[4]));
  AL_DFF_X al_31f2bc3d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c8474427[5]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_8c490204[5]));
  AL_DFF_X al_5c576f1f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c8474427[6]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_8c490204[6]));
  AL_DFF_X al_53496a4b (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c8474427[7]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_8c490204[7]));
  AL_DFF_X al_413d5334 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c8474427[8]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_8c490204[8]));
  AL_DFF_X al_8d8da18e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_63a836a9[0]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_24ac8493[0]));
  AL_DFF_X al_f13f0dd7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_63a836a9[1]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_24ac8493[1]));
  AL_DFF_X al_af5588d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_63a836a9[2]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_24ac8493[2]));
  AL_DFF_X al_a9378f0a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c122424e[0]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_54d2aa3[0]));
  AL_DFF_X al_638e8f14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c122424e[1]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_54d2aa3[1]));
  AL_DFF_X al_c772c33c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c122424e[2]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_54d2aa3[2]));
  AL_DFF_X al_545c3cf7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c122424e[3]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_54d2aa3[3]));
  AL_DFF_X al_e2ab8394 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c122424e[4]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_54d2aa3[4]));
  AL_DFF_X al_aceaebac (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c122424e[5]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_54d2aa3[5]));
  AL_DFF_X al_893deeb5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c122424e[6]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_54d2aa3[6]));
  AL_DFF_X al_1952da23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c122424e[7]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_54d2aa3[7]));
  AL_DFF_X al_eaa51de5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b3968bab[0]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_77f0ddfc[0]));
  AL_DFF_X al_4849d172 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_b3968bab[1]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_77f0ddfc[1]));
  AL_DFF_X al_8245c217 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_630a3426[0]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_f3f63e4d[0]));
  AL_DFF_X al_7575b1ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_630a3426[1]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_f3f63e4d[1]));
  AL_DFF_X al_a19ad63d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_77695f5b[0]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_e8bb9040[0]));
  AL_DFF_X al_baaafe79 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_77695f5b[9]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_e8bb9040[9]));
  AL_DFF_X al_3b50f921 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_77695f5b[10]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_e8bb9040[10]));
  AL_DFF_X al_cd41d57e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_77695f5b[11]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_e8bb9040[11]));
  AL_DFF_X al_33424807 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_77695f5b[12]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_e8bb9040[12]));
  AL_DFF_X al_e7bd4dcb (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_77695f5b[13]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_e8bb9040[13]));
  AL_DFF_X al_f37ed438 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_77695f5b[14]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_e8bb9040[14]));
  AL_DFF_X al_c655741a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_77695f5b[15]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_e8bb9040[15]));
  AL_DFF_X al_aad72f5d (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_77695f5b[16]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_e8bb9040[16]));
  AL_DFF_X al_c3e18a5a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_77695f5b[17]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_e8bb9040[17]));
  AL_DFF_X al_64a3ee71 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_77695f5b[18]),
    .en(tx_clk_en),
    .sr(al_6b4499fc),
    .ss(1'b0),
    .q(al_e8bb9040[18]));
  AL_DFF_X al_f0ed4056 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_77695f5b[1]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_e8bb9040[1]));
  AL_DFF_X al_fccb2998 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_77695f5b[2]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_e8bb9040[2]));
  AL_DFF_X al_63773dbe (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_77695f5b[3]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_e8bb9040[3]));
  AL_DFF_X al_a83e820f (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_77695f5b[4]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_e8bb9040[4]));
  AL_DFF_X al_2c70d3eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_77695f5b[5]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_e8bb9040[5]));
  AL_DFF_X al_86f41d7e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_77695f5b[6]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_e8bb9040[6]));
  AL_DFF_X al_565c9074 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_77695f5b[7]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_e8bb9040[7]));
  AL_DFF_X al_d318fb15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_77695f5b[8]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_e8bb9040[8]));
  AL_DFF_X al_2c129b43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_20b55994[0]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_5f257019[0]));
  AL_DFF_X al_36dcf325 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_20b55994[1]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_5f257019[1]));
  AL_DFF_X al_5703b70e (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_20b55994[2]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_5f257019[2]));
  AL_DFF_X al_e00fdec6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_20b55994[3]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_5f257019[3]));
  AL_DFF_X al_efe8e24c (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_20b55994[4]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_5f257019[4]));
  AL_DFF_X al_1d422ad7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_20b55994[5]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(al_6b4499fc),
    .q(al_5f257019[5]));
  AL_DFF_X al_1b16ca13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c007c6a1[0]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e512aff[0]));
  AL_DFF_X al_19c97f36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c007c6a1[9]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e512aff[9]));
  AL_DFF_X al_82cf3fcd (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c007c6a1[10]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e512aff[10]));
  AL_DFF_X al_ecaa6e15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c007c6a1[11]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e512aff[11]));
  AL_DFF_X al_fa471567 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c007c6a1[12]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e512aff[12]));
  AL_DFF_X al_e030ac3a (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c007c6a1[13]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e512aff[13]));
  AL_DFF_X al_8ead11f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c007c6a1[14]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e512aff[14]));
  AL_DFF_X al_c00d14e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c007c6a1[1]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e512aff[1]));
  AL_DFF_X al_a09d44ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c007c6a1[2]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e512aff[2]));
  AL_DFF_X al_6833a615 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c007c6a1[3]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e512aff[3]));
  AL_DFF_X al_ec59eca7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c007c6a1[4]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e512aff[4]));
  AL_DFF_X al_58a4a279 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c007c6a1[5]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e512aff[5]));
  AL_DFF_X al_cb886a26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c007c6a1[6]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e512aff[6]));
  AL_DFF_X al_1fb87d18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c007c6a1[7]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e512aff[7]));
  AL_DFF_X al_a66180b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(tx_mac_clk),
    .d(al_c007c6a1[8]),
    .en(tx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e512aff[8]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_9799382b (
    .a(1'b0),
    .o({al_7868fcca,open_n18}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a6cc7cef (
    .a(al_e8bb9040[0]),
    .b(1'b1),
    .c(al_7868fcca),
    .o({al_78567007,al_acbf9207[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f6900725 (
    .a(al_e8bb9040[1]),
    .b(1'b0),
    .c(al_78567007),
    .o({al_3efdaf7e,al_acbf9207[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1b408c6b (
    .a(al_e8bb9040[2]),
    .b(1'b0),
    .c(al_3efdaf7e),
    .o({al_e4a226df,al_acbf9207[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c6e4f315 (
    .a(al_e8bb9040[3]),
    .b(1'b0),
    .c(al_e4a226df),
    .o({al_dbdccc1f,al_acbf9207[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4722be8d (
    .a(al_e8bb9040[4]),
    .b(1'b0),
    .c(al_dbdccc1f),
    .o({al_9bcb8f17,al_acbf9207[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_db937b4a (
    .a(al_e8bb9040[5]),
    .b(1'b0),
    .c(al_9bcb8f17),
    .o({al_81191a79,al_acbf9207[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_59c93334 (
    .a(al_e8bb9040[6]),
    .b(1'b0),
    .c(al_81191a79),
    .o({al_a6edfc2,al_acbf9207[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bfa3b596 (
    .a(al_e8bb9040[7]),
    .b(1'b0),
    .c(al_a6edfc2),
    .o({al_3abe5c64,al_acbf9207[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cd2e9eb5 (
    .a(al_e8bb9040[8]),
    .b(1'b0),
    .c(al_3abe5c64),
    .o({al_f974815d,al_acbf9207[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_379c4bbc (
    .a(al_e8bb9040[9]),
    .b(1'b0),
    .c(al_f974815d),
    .o({al_7f233c39,al_acbf9207[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4785fc74 (
    .a(al_e8bb9040[10]),
    .b(1'b0),
    .c(al_7f233c39),
    .o({al_42136331,al_acbf9207[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_355c869b (
    .a(al_e8bb9040[11]),
    .b(1'b0),
    .c(al_42136331),
    .o({al_5832a18a,al_acbf9207[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1e7507c9 (
    .a(al_e8bb9040[12]),
    .b(1'b0),
    .c(al_5832a18a),
    .o({al_fde4e9e1,al_acbf9207[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7bb3740e (
    .a(al_e8bb9040[13]),
    .b(1'b0),
    .c(al_fde4e9e1),
    .o({al_6b963607,al_acbf9207[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3be1eb48 (
    .a(al_e8bb9040[14]),
    .b(1'b0),
    .c(al_6b963607),
    .o({al_e364ec9e,al_acbf9207[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3231a0bc (
    .a(al_e8bb9040[15]),
    .b(1'b0),
    .c(al_e364ec9e),
    .o({al_923f48aa,al_acbf9207[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_68558a0a (
    .a(al_e8bb9040[16]),
    .b(1'b0),
    .c(al_923f48aa),
    .o({al_7b831e20,al_acbf9207[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8fc658e (
    .a(al_e8bb9040[17]),
    .b(1'b0),
    .c(al_7b831e20),
    .o({al_4d9c1d5,al_acbf9207[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f75581c8 (
    .a(al_e8bb9040[18]),
    .b(1'b0),
    .c(al_4d9c1d5),
    .o({open_n19,al_acbf9207[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_6d220656 (
    .a(1'b0),
    .o({al_ec490bfd,open_n22}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9a8a00eb (
    .a(al_8e462c61[0]),
    .b(1'b1),
    .c(al_ec490bfd),
    .o({al_58bd59f6,al_e20fd0c7[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b0300ffb (
    .a(al_8e462c61[1]),
    .b(1'b0),
    .c(al_58bd59f6),
    .o({al_ebd456eb,al_e20fd0c7[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cb3e4530 (
    .a(al_8e462c61[2]),
    .b(1'b0),
    .c(al_ebd456eb),
    .o({al_b59c2e50,al_e20fd0c7[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_26107a32 (
    .a(al_8e462c61[3]),
    .b(1'b0),
    .c(al_b59c2e50),
    .o({al_575bbbae,al_e20fd0c7[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_50551443 (
    .a(al_8e462c61[4]),
    .b(1'b0),
    .c(al_575bbbae),
    .o({al_6f9895cd,al_e20fd0c7[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_225abe (
    .a(al_8e462c61[5]),
    .b(1'b0),
    .c(al_6f9895cd),
    .o({al_b0d2bfc8,al_e20fd0c7[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6746cc98 (
    .a(al_8e462c61[6]),
    .b(1'b0),
    .c(al_b0d2bfc8),
    .o({al_73782b81,al_e20fd0c7[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_335cf46b (
    .a(al_8e462c61[7]),
    .b(1'b0),
    .c(al_73782b81),
    .o({al_29cb65c6,al_e20fd0c7[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cc1dfa54 (
    .a(al_8e462c61[8]),
    .b(1'b0),
    .c(al_29cb65c6),
    .o({al_7a2a1104,al_e20fd0c7[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3120ca90 (
    .a(al_8e462c61[9]),
    .b(1'b0),
    .c(al_7a2a1104),
    .o({al_1e9fbff4,al_e20fd0c7[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5a1baede (
    .a(al_8e462c61[10]),
    .b(1'b0),
    .c(al_1e9fbff4),
    .o({al_d2811bd8,al_e20fd0c7[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_58b252b3 (
    .a(al_8e462c61[11]),
    .b(1'b0),
    .c(al_d2811bd8),
    .o({al_f2cdbc14,al_e20fd0c7[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bc21601b (
    .a(al_8e462c61[12]),
    .b(1'b0),
    .c(al_f2cdbc14),
    .o({al_fc353ce9,al_e20fd0c7[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9c8499fa (
    .a(al_8e462c61[13]),
    .b(1'b0),
    .c(al_fc353ce9),
    .o({al_dfffc03a,al_e20fd0c7[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6abf855e (
    .a(al_8e462c61[14]),
    .b(1'b0),
    .c(al_dfffc03a),
    .o({open_n23,al_e20fd0c7[14]}));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_bbf8458 (
    .a(al_b984f6c1),
    .b(al_9b4eaefc[4]),
    .o(al_fadd6423));
  AL_DFF_X al_9ebd276 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_114295f1),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_4596a396));
  AL_DFF_X al_6ed82bec (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1c6db97d),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_dbe2baa6));
  AL_DFF_X al_37753f90 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_56997d45),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_7bec6b72));
  AL_DFF_X al_d5042958 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_132ae268),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_30b5e311));
  AL_DFF_0 al_bfa93eb5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_59a83809),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ecfcb422[0]));
  AL_DFF_0 al_70af7f40 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ecfcb422[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ecfcb422[1]));
  AL_DFF_0 al_70d83c24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ecfcb422[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ecfcb422[2]));
  AL_DFF_0 al_ead9b1d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ecfcb422[2]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ecfcb422[3]));
  AL_DFF_X al_65033afe (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_e4f9c44c),
    .en(1'b1),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_a9336f5));
  AL_DFF_X al_59b8947d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1430ac7c),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f15a934));
  AL_DFF_X al_a36db9a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f452d0ae),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b5e36a9));
  AL_DFF_X al_a0342538 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_33c6f6),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d976dda9));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*B*A)"),
    .INIT(64'h0000000000000008))
    al_1a8358c (
    .a(al_5ec57682),
    .b(al_41ffdcd4),
    .c(al_13660933[0]),
    .d(al_13660933[1]),
    .e(al_13660933[4]),
    .f(al_13660933[5]),
    .o(al_78991444));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*~B*A)"),
    .INIT(32'h00000020))
    al_922f0546 (
    .a(al_78991444),
    .b(al_b9297703[0]),
    .c(al_b9297703[1]),
    .d(al_b9297703[2]),
    .e(al_b9297703[3]),
    .o(al_8f82c712));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    al_47c42dc0 (
    .a(al_78991444),
    .b(al_b9297703[0]),
    .c(al_b9297703[1]),
    .d(al_b9297703[2]),
    .e(al_b9297703[3]),
    .o(al_82faa065));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    al_ace91a7b (
    .a(al_78991444),
    .b(al_b9297703[0]),
    .c(al_b9297703[1]),
    .d(al_b9297703[2]),
    .e(al_b9297703[3]),
    .o(al_b7164eee));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    al_fea4ebab (
    .a(al_134c8dab),
    .b(al_b9297703[0]),
    .c(al_b9297703[1]),
    .d(al_b9297703[2]),
    .e(al_b9297703[3]),
    .o(al_e3838f69));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    al_1b2c3158 (
    .a(al_134c8dab),
    .b(al_b9297703[0]),
    .c(al_b9297703[1]),
    .d(al_b9297703[2]),
    .e(al_b9297703[3]),
    .o(al_4965e5fa));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_2d618b87 (
    .a(s_axi_awvalid),
    .b(s_axi_wvalid),
    .c(s_axi_wready),
    .o(al_5df5c44f));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_ad3f31fd (
    .a(al_13660933[6]),
    .b(al_13660933[7]),
    .o(al_41ffdcd4));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*~B*A)"),
    .INIT(32'h00000020))
    al_e92faa67 (
    .a(al_41ffdcd4),
    .b(al_13660933[0]),
    .c(al_13660933[1]),
    .d(al_13660933[4]),
    .e(al_13660933[5]),
    .o(al_7afe69f4));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~B*A*~(D*C))"),
    .INIT(64'h0000000000000222))
    al_4be83be3 (
    .a(al_13660933[2]),
    .b(al_13660933[3]),
    .c(al_b9297703[0]),
    .d(al_b9297703[1]),
    .e(al_b9297703[2]),
    .f(al_b9297703[3]),
    .o(al_74a15ab1));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_5c758555 (
    .a(al_74a15ab1),
    .b(al_5df5c44f),
    .o(al_5ec57682));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_34f2fff1 (
    .a(al_5ec57682),
    .b(al_7afe69f4),
    .o(al_134c8dab));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*~B*A)"),
    .INIT(32'h00000020))
    al_c5940a5a (
    .a(al_134c8dab),
    .b(al_b9297703[0]),
    .c(al_b9297703[1]),
    .d(al_b9297703[2]),
    .e(al_b9297703[3]),
    .o(al_71f17e1a));
  AL_MAP_LUT6 #(
    .EQN("((D*~(F)*~((C*B))+D*F*~((C*B))+~(D)*F*(C*B)+D*F*(C*B))*~(~E*A))"),
    .INIT(64'hffc055403f001500))
    al_21fb12be (
    .a(al_132ae268),
    .b(al_968fd17c),
    .c(al_d0555e9d[2]),
    .d(al_8399b753),
    .e(al_30b5e311),
    .f(al_3edda74b),
    .o(al_1bc55ab2));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    al_115bd025 (
    .a(al_a03de72f),
    .b(al_88fb5330[16]),
    .c(al_a9336f5),
    .o(al_e6b493f[16]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    al_eca98982 (
    .a(al_81681eb),
    .b(al_88fb5330[17]),
    .c(al_a9336f5),
    .o(al_e6b493f[17]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    al_94a79df8 (
    .a(al_644f021d),
    .b(al_88fb5330[18]),
    .c(al_a9336f5),
    .o(al_e6b493f[18]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    al_b177a56e (
    .a(al_f4252f15),
    .b(al_88fb5330[19]),
    .c(al_a9336f5),
    .o(al_e6b493f[19]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    al_b047ea29 (
    .a(al_61fb0a6),
    .b(al_88fb5330[20]),
    .c(al_a9336f5),
    .o(al_e6b493f[20]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    al_d5ce5d81 (
    .a(al_3b505c23),
    .b(al_88fb5330[21]),
    .c(al_a9336f5),
    .o(al_e6b493f[21]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    al_a23c580 (
    .a(al_179835d0),
    .b(al_88fb5330[22]),
    .c(al_a9336f5),
    .o(al_e6b493f[22]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    al_4054bb78 (
    .a(al_7cd2fee3),
    .b(al_88fb5330[23]),
    .c(al_a9336f5),
    .o(al_e6b493f[23]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    al_d25f08e4 (
    .a(al_70727c2f),
    .b(al_88fb5330[24]),
    .c(al_a9336f5),
    .o(al_e6b493f[24]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    al_f8eee492 (
    .a(al_e5314cad),
    .b(al_88fb5330[25]),
    .c(al_a9336f5),
    .o(al_e6b493f[25]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    al_50543807 (
    .a(al_70372a24),
    .b(al_88fb5330[26]),
    .c(al_a9336f5),
    .o(al_e6b493f[26]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    al_581d58bb (
    .a(al_1824196b),
    .b(al_88fb5330[27]),
    .c(al_a9336f5),
    .o(al_e6b493f[27]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    al_1ac8a80 (
    .a(al_67074a64),
    .b(al_88fb5330[28]),
    .c(al_a9336f5),
    .o(al_e6b493f[28]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    al_e5ccd36e (
    .a(al_737a8715),
    .b(al_88fb5330[29]),
    .c(al_a9336f5),
    .o(al_e6b493f[29]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    al_84f8c05c (
    .a(al_90021ccb),
    .b(al_88fb5330[30]),
    .c(al_a9336f5),
    .o(al_e6b493f[30]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    al_ead443c7 (
    .a(al_4c4d90b0),
    .b(al_88fb5330[31]),
    .c(al_a9336f5),
    .o(al_e6b493f[31]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_576e007e (
    .a(al_7bce675b),
    .b(al_9e8909aa),
    .o(al_132ae268));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F)"),
    .INIT(64'h32f336f73afb3eff))
    al_dee712d7 (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_d0555e9d[2]),
    .d(al_752f7592[7]),
    .e(al_752f7592[23]),
    .f(al_752f7592[31]),
    .o(al_8ab6e600));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_7787b3d8 (
    .a(al_d0555e9d[0]),
    .b(al_752f7592[36]),
    .c(al_752f7592[44]),
    .o(al_4974667d));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_fdf4ae7 (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_752f7592[4]),
    .d(al_752f7592[12]),
    .e(al_752f7592[20]),
    .f(al_752f7592[28]),
    .o(al_3255583f));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff3fafaf0030a0a0))
    al_5298bf68 (
    .a(al_3255583f),
    .b(al_4974667d),
    .c(al_132ae268),
    .d(al_d0555e9d[1]),
    .e(al_d0555e9d[2]),
    .f(al_752f7592[4]),
    .o(al_3a736cff[4]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_783d1ab (
    .a(al_d0555e9d[0]),
    .b(al_752f7592[37]),
    .c(al_752f7592[45]),
    .o(al_fd84e521));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_9357c9fd (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_752f7592[5]),
    .d(al_752f7592[13]),
    .e(al_752f7592[21]),
    .f(al_752f7592[29]),
    .o(al_b91e0498));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff3fafaf0030a0a0))
    al_50f06a13 (
    .a(al_b91e0498),
    .b(al_fd84e521),
    .c(al_132ae268),
    .d(al_d0555e9d[1]),
    .e(al_d0555e9d[2]),
    .f(al_752f7592[5]),
    .o(al_3a736cff[5]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_3f05a2d1 (
    .a(al_132ae268),
    .b(al_d0555e9d[0]),
    .c(al_d0555e9d[1]),
    .d(al_d0555e9d[2]),
    .o(al_9b5719ae));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_d01a99dd (
    .a(al_d0555e9d[0]),
    .b(al_752f7592[34]),
    .c(al_752f7592[42]),
    .o(al_1f5e6438));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_e9a7124d (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_752f7592[2]),
    .d(al_752f7592[10]),
    .e(al_752f7592[18]),
    .f(al_752f7592[26]),
    .o(al_67edee18));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff3fafaf0030a0a0))
    al_9f8b70a2 (
    .a(al_67edee18),
    .b(al_1f5e6438),
    .c(al_132ae268),
    .d(al_d0555e9d[1]),
    .e(al_d0555e9d[2]),
    .f(al_752f7592[2]),
    .o(al_3a736cff[2]));
  AL_MAP_LUT6 #(
    .EQN("(~B*(A*~(C)*D*~(E)*~(F)+~(A)*C*~(D)*E*~(F)+A*~(C)*D*E*~(F)+~(A)*C*D*E*~(F)+A*C*~(D)*~(E)*F+A*~(C)*D*~(E)*F+A*C*D*~(E)*F+~(A)*C*~(D)*E*F+A*C*~(D)*E*F+A*~(C)*D*E*F+~(A)*C*D*E*F+A*C*D*E*F))"),
    .INIT(64'h3230222012100200))
    al_1f85d042 (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_d0555e9d[2]),
    .d(al_752f7592[14]),
    .e(al_752f7592[38]),
    .f(al_752f7592[46]),
    .o(al_e410470b));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F)"),
    .INIT(64'h32f336f73afb3eff))
    al_778a9553 (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_d0555e9d[2]),
    .d(al_752f7592[6]),
    .e(al_752f7592[22]),
    .f(al_752f7592[30]),
    .o(al_587ea99f));
  AL_MAP_LUT6 #(
    .EQN("(~B*(A*~(C)*D*~(E)*~(F)+~(A)*C*~(D)*E*~(F)+A*~(C)*D*E*~(F)+~(A)*C*D*E*~(F)+A*C*~(D)*~(E)*F+A*~(C)*D*~(E)*F+A*C*D*~(E)*F+~(A)*C*~(D)*E*F+A*C*~(D)*E*F+A*~(C)*D*E*F+~(A)*C*D*E*F+A*C*D*E*F))"),
    .INIT(64'h3230222012100200))
    al_3beca40 (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_d0555e9d[2]),
    .d(al_752f7592[11]),
    .e(al_752f7592[35]),
    .f(al_752f7592[43]),
    .o(al_6bff803e));
  AL_MAP_LUT5 #(
    .EQN("(~C*B*(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))"),
    .INIT(32'h0c080400))
    al_21f15610 (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_d0555e9d[2]),
    .d(al_752f7592[19]),
    .e(al_752f7592[27]),
    .o(al_2a3de543));
  AL_MAP_LUT5 #(
    .EQN("(E*~(A*(B*~(C)*~(D)+~(B)*C*~(D)+B*C*~(D)+~(B)*~(C)*D+B*~(C)*D)))"),
    .INIT(32'hf5570000))
    al_53fce6a6 (
    .a(al_132ae268),
    .b(al_d0555e9d[0]),
    .c(al_d0555e9d[1]),
    .d(al_d0555e9d[2]),
    .e(al_752f7592[3]),
    .o(al_5716efe6));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_3d31b267 (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_752f7592[0]),
    .d(al_752f7592[8]),
    .e(al_752f7592[16]),
    .f(al_752f7592[24]),
    .o(al_d9e64745));
  AL_MAP_LUT6 #(
    .EQN("~(A*~((~C*(E*~(F)*~(B)+E*F*~(B)+~(E)*F*B+E*F*B)))*~(D)+A*(~C*(E*~(F)*~(B)+E*F*~(B)+~(E)*F*B+E*F*B))*~(D)+~(A)*(~C*(E*~(F)*~(B)+E*F*~(B)+~(E)*F*B+E*F*B))*D+A*(~C*(E*~(F)*~(B)+E*F*~(B)+~(E)*F*B+E*F*B))*D)"),
    .INIT(64'hf055f355fc55ff55))
    al_7bf102ee (
    .a(al_d9e64745),
    .b(al_d0555e9d[0]),
    .c(al_d0555e9d[1]),
    .d(al_d0555e9d[2]),
    .e(al_752f7592[32]),
    .f(al_752f7592[40]),
    .o(al_70d272c9));
  AL_MAP_LUT5 #(
    .EQN("~(E@(~A*~(D*~(~C*~B))))"),
    .INIT(32'h0155feaa))
    al_1b231817 (
    .a(al_5716efe6),
    .b(al_6bff803e),
    .c(al_2a3de543),
    .d(al_132ae268),
    .e(al_e8c5f626[3]),
    .o(al_b17db8f));
  AL_MAP_LUT6 #(
    .EQN("(C@(~(A)*B*~((E*D))*~(F)+~(A)*B*(E*D)*~(F)+~(A)*~(B)*~((E*D))*F+A*~(B)*~((E*D))*F+~(A)*B*~((E*D))*F+~(A)*~(B)*(E*D)*F+A*~(B)*(E*D)*F+~(A)*B*(E*D)*F+A*B*(E*D)*F))"),
    .INIT(64'h0f878787b4b4b4b4))
    al_bdb66821 (
    .a(al_70d272c9),
    .b(al_132ae268),
    .c(al_e8c5f626[0]),
    .d(al_d0555e9d[1]),
    .e(al_d0555e9d[2]),
    .f(al_752f7592[0]),
    .o(al_740a6bb3));
  AL_MAP_LUT5 #(
    .EQN("(D@(~E*~((B*~A))*~(C)+~E*(B*~A)*~(C)+~(~E)*(B*~A)*C+~E*(B*~A)*C))"),
    .INIT(32'hbf40b04f))
    al_d2c0145a (
    .a(al_e410470b),
    .b(al_587ea99f),
    .c(al_132ae268),
    .d(al_e8c5f626[6]),
    .e(al_752f7592[6]),
    .o(al_7b32ad34));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_bd88ed58 (
    .a(al_d0555e9d[0]),
    .b(al_752f7592[33]),
    .c(al_752f7592[41]),
    .o(al_f2d1cf9));
  AL_MAP_LUT6 #(
    .EQN("(~(E@C)*~(F@B)*~(D@A))"),
    .INIT(64'h8040080420100201))
    al_699b40f5 (
    .a(al_3a736cff[1]),
    .b(al_3a736cff[4]),
    .c(al_3a736cff[2]),
    .d(al_e8c5f626[1]),
    .e(al_e8c5f626[2]),
    .f(al_e8c5f626[4]),
    .o(al_ab134353));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B@A))"),
    .INIT(8'h90))
    al_ad587093 (
    .a(al_3a736cff[5]),
    .b(al_e8c5f626[5]),
    .c(al_8f15a934),
    .o(al_3eaa9cdd));
  AL_MAP_LUT6 #(
    .EQN("(A*(E@(~F*~((C*~B))*~(D)+~F*(C*~B)*~(D)+~(~F)*(C*~B)*D+~F*(C*~B)*D)))"),
    .INIT(64'h8aaa20008a0020aa))
    al_a2f697d5 (
    .a(al_7b32ad34),
    .b(al_7be18307),
    .c(al_8ab6e600),
    .d(al_132ae268),
    .e(al_e8c5f626[7]),
    .f(al_752f7592[7]),
    .o(al_53669626));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(~E*D*~C*B*A))"),
    .INIT(64'hffffffff00000800))
    al_6cc0eabf (
    .a(al_ab134353),
    .b(al_53669626),
    .c(al_740a6bb3),
    .d(al_3eaa9cdd),
    .e(al_b17db8f),
    .f(al_9b5719ae),
    .o(al_1430ac7c));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_16b2aa3c (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_752f7592[1]),
    .d(al_752f7592[9]),
    .e(al_752f7592[17]),
    .f(al_752f7592[25]),
    .o(al_47ed325a));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff3fafaf0030a0a0))
    al_62d599f (
    .a(al_47ed325a),
    .b(al_f2d1cf9),
    .c(al_132ae268),
    .d(al_d0555e9d[1]),
    .e(al_d0555e9d[2]),
    .f(al_752f7592[1]),
    .o(al_3a736cff[1]));
  AL_MAP_LUT6 #(
    .EQN("(~B*(A*~(C)*D*~(E)*~(F)+~(A)*C*~(D)*E*~(F)+A*~(C)*D*E*~(F)+~(A)*C*D*E*~(F)+A*C*~(D)*~(E)*F+A*~(C)*D*~(E)*F+A*C*D*~(E)*F+~(A)*C*~(D)*E*F+A*C*~(D)*E*F+A*~(C)*D*E*F+~(A)*C*D*E*F+A*C*D*E*F))"),
    .INIT(64'h3230222012100200))
    al_ff286764 (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_d0555e9d[2]),
    .d(al_752f7592[15]),
    .e(al_752f7592[39]),
    .f(al_752f7592[47]),
    .o(al_7be18307));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_32336675 (
    .a(al_d0555e9d[0]),
    .b(al_d1b76c6b[34]),
    .c(al_d1b76c6b[42]),
    .o(al_edebc70b));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F)"),
    .INIT(64'h32f336f73afb3eff))
    al_a97f428c (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_d0555e9d[2]),
    .d(al_d1b76c6b[6]),
    .e(al_d1b76c6b[22]),
    .f(al_d1b76c6b[30]),
    .o(al_8d4887c7));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_12c31040 (
    .a(al_d0555e9d[0]),
    .b(al_d1b76c6b[37]),
    .c(al_d1b76c6b[45]),
    .o(al_aaacabd5));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_2cff8143 (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_d1b76c6b[5]),
    .d(al_d1b76c6b[13]),
    .e(al_d1b76c6b[21]),
    .f(al_d1b76c6b[29]),
    .o(al_c7b03fcb));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff3fafaf0030a0a0))
    al_fea6d7b (
    .a(al_c7b03fcb),
    .b(al_aaacabd5),
    .c(al_132ae268),
    .d(al_d0555e9d[1]),
    .e(al_d0555e9d[2]),
    .f(al_d1b76c6b[5]),
    .o(al_3a736cff[13]));
  AL_MAP_LUT6 #(
    .EQN("(~B*(A*~(C)*D*~(E)*~(F)+~(A)*C*~(D)*E*~(F)+A*~(C)*D*E*~(F)+~(A)*C*D*E*~(F)+A*C*~(D)*~(E)*F+A*~(C)*D*~(E)*F+A*C*D*~(E)*F+~(A)*C*~(D)*E*F+A*C*~(D)*E*F+A*~(C)*D*E*F+~(A)*C*D*E*F+A*C*D*E*F))"),
    .INIT(64'h3230222012100200))
    al_72637ff3 (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_d0555e9d[2]),
    .d(al_d1b76c6b[11]),
    .e(al_d1b76c6b[35]),
    .f(al_d1b76c6b[43]),
    .o(al_1ec4cd29));
  AL_MAP_LUT5 #(
    .EQN("(~C*B*(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))"),
    .INIT(32'h0c080400))
    al_a41a7b16 (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_d0555e9d[2]),
    .d(al_d1b76c6b[19]),
    .e(al_d1b76c6b[27]),
    .o(al_88a2bdf0));
  AL_MAP_LUT5 #(
    .EQN("(E*~(A*(B*~(C)*~(D)+~(B)*C*~(D)+B*C*~(D)+~(B)*~(C)*D+B*~(C)*D)))"),
    .INIT(32'hf5570000))
    al_7895e38 (
    .a(al_132ae268),
    .b(al_d0555e9d[0]),
    .c(al_d0555e9d[1]),
    .d(al_d0555e9d[2]),
    .e(al_d1b76c6b[3]),
    .o(al_468d7712));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_308dbbee (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_d1b76c6b[0]),
    .d(al_d1b76c6b[8]),
    .e(al_d1b76c6b[16]),
    .f(al_d1b76c6b[24]),
    .o(al_ec16c3b2));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_b1d7c8c1 (
    .a(al_d0555e9d[0]),
    .b(al_d1b76c6b[32]),
    .c(al_d1b76c6b[40]),
    .o(al_1b37ba12));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00c05050ffcf5f5f))
    al_a31d9dd7 (
    .a(al_ec16c3b2),
    .b(al_1b37ba12),
    .c(al_132ae268),
    .d(al_d0555e9d[1]),
    .e(al_d0555e9d[2]),
    .f(al_d1b76c6b[0]),
    .o(al_9c1262a5));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    al_46931b6b (
    .a(al_9c1262a5),
    .b(al_e8c5f626[0]),
    .o(al_fcec21f3));
  AL_MAP_LUT6 #(
    .EQN("(~B*(A*~(C)*D*~(E)*~(F)+~(A)*C*~(D)*E*~(F)+A*~(C)*D*E*~(F)+~(A)*C*D*E*~(F)+A*C*~(D)*~(E)*F+A*~(C)*D*~(E)*F+A*C*D*~(E)*F+~(A)*C*~(D)*E*F+A*C*~(D)*E*F+A*~(C)*D*E*F+~(A)*C*D*E*F+A*C*D*E*F))"),
    .INIT(64'h3230222012100200))
    al_5335f2b (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_d0555e9d[2]),
    .d(al_d1b76c6b[15]),
    .e(al_d1b76c6b[39]),
    .f(al_d1b76c6b[47]),
    .o(al_39bb30c0));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_10191a75 (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_d1b76c6b[2]),
    .d(al_d1b76c6b[10]),
    .e(al_d1b76c6b[18]),
    .f(al_d1b76c6b[26]),
    .o(al_65907c46));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F)"),
    .INIT(64'h32f336f73afb3eff))
    al_4ee3a952 (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_d0555e9d[2]),
    .d(al_d1b76c6b[7]),
    .e(al_d1b76c6b[23]),
    .f(al_d1b76c6b[31]),
    .o(al_d6e69fcf));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_f69a67dd (
    .a(al_d0555e9d[0]),
    .b(al_d1b76c6b[36]),
    .c(al_d1b76c6b[44]),
    .o(al_3b01668f));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_3f461560 (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_d1b76c6b[4]),
    .d(al_d1b76c6b[12]),
    .e(al_d1b76c6b[20]),
    .f(al_d1b76c6b[28]),
    .o(al_5c5a5e75));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff3fafaf0030a0a0))
    al_9e4670f2 (
    .a(al_5c5a5e75),
    .b(al_3b01668f),
    .c(al_132ae268),
    .d(al_d0555e9d[1]),
    .e(al_d0555e9d[2]),
    .f(al_d1b76c6b[4]),
    .o(al_3a736cff[12]));
  AL_MAP_LUT5 #(
    .EQN("~(E@(~A*~(D*~(~C*~B))))"),
    .INIT(32'h0155feaa))
    al_94917954 (
    .a(al_468d7712),
    .b(al_1ec4cd29),
    .c(al_88a2bdf0),
    .d(al_132ae268),
    .e(al_e8c5f626[3]),
    .o(al_8e2b6222));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    al_9da0dc4e (
    .a(al_3a736cff[13]),
    .b(al_e8c5f626[5]),
    .o(al_1e78f688));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff3fafaf0030a0a0))
    al_fcfd284b (
    .a(al_65907c46),
    .b(al_edebc70b),
    .c(al_132ae268),
    .d(al_d0555e9d[1]),
    .e(al_d0555e9d[2]),
    .f(al_d1b76c6b[2]),
    .o(al_3a736cff[10]));
  AL_MAP_LUT6 #(
    .EQN("(F*~B*~(E@C)*~(D@A))"),
    .INIT(64'h2010020100000000))
    al_39c5fae9 (
    .a(al_3a736cff[10]),
    .b(al_b1b43431),
    .c(al_3a736cff[12]),
    .d(al_e8c5f626[2]),
    .e(al_e8c5f626[4]),
    .f(al_b5e36a9),
    .o(al_13600bf4));
  AL_MAP_LUT5 #(
    .EQN("(D@(~E*~((B*~A))*~(C)+~E*(B*~A)*~(C)+~(~E)*(B*~A)*C+~E*(B*~A)*C))"),
    .INIT(32'hbf40b04f))
    al_4723062d (
    .a(al_39bb30c0),
    .b(al_d6e69fcf),
    .c(al_132ae268),
    .d(al_e8c5f626[7]),
    .e(al_d1b76c6b[7]),
    .o(al_5bb5921));
  AL_MAP_LUT6 #(
    .EQN("(A*(E@(~F*~((C*~B))*~(D)+~F*(C*~B)*~(D)+~(~F)*(C*~B)*D+~F*(C*~B)*D)))"),
    .INIT(64'h8aaa20008a0020aa))
    al_6788ae3c (
    .a(al_5bb5921),
    .b(al_e6700530),
    .c(al_8d4887c7),
    .d(al_132ae268),
    .e(al_e8c5f626[6]),
    .f(al_d1b76c6b[6]),
    .o(al_a024e6ee));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(~E*D*C*B*A))"),
    .INIT(64'hffffffff00008000))
    al_5cfa163d (
    .a(al_13600bf4),
    .b(al_a024e6ee),
    .c(al_fcec21f3),
    .d(al_1e78f688),
    .e(al_8e2b6222),
    .f(al_9b5719ae),
    .o(al_f452d0ae));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*~(C)*~(B)+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*~(B)+~((D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))*C*B+(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A)*C*B)"),
    .INIT(32'hf3e2d1c0))
    al_b8d6b9c7 (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_d1b76c6b[1]),
    .d(al_d1b76c6b[33]),
    .e(al_d1b76c6b[41]),
    .o(al_2f3d50c1));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_c4ade397 (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_d1b76c6b[1]),
    .d(al_d1b76c6b[9]),
    .e(al_d1b76c6b[17]),
    .f(al_d1b76c6b[25]),
    .o(al_71c12aaa));
  AL_MAP_LUT6 #(
    .EQN("(D@(F*~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*~(C)+F*(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)+~(F)*(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C+F*(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C))"),
    .INIT(64'h30cf50af3fc05fa0))
    al_bf9961d6 (
    .a(al_71c12aaa),
    .b(al_2f3d50c1),
    .c(al_132ae268),
    .d(al_e8c5f626[1]),
    .e(al_d0555e9d[2]),
    .f(al_d1b76c6b[1]),
    .o(al_b1b43431));
  AL_MAP_LUT6 #(
    .EQN("(~B*(A*~(C)*D*~(E)*~(F)+~(A)*C*~(D)*E*~(F)+A*~(C)*D*E*~(F)+~(A)*C*D*E*~(F)+A*C*~(D)*~(E)*F+A*~(C)*D*~(E)*F+A*C*D*~(E)*F+~(A)*C*~(D)*E*F+A*C*~(D)*E*F+A*~(C)*D*E*F+~(A)*C*D*E*F+A*C*D*E*F))"),
    .INIT(64'h3230222012100200))
    al_552ff953 (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_d0555e9d[2]),
    .d(al_d1b76c6b[14]),
    .e(al_d1b76c6b[38]),
    .f(al_d1b76c6b[46]),
    .o(al_e6700530));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_5164e042 (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_902efd00[6]),
    .d(al_902efd00[14]),
    .e(al_902efd00[22]),
    .f(al_902efd00[30]),
    .o(al_2cc28140));
  AL_MAP_LUT5 #(
    .EQN("~(E@(~B*~(D*~(~C*~A))))"),
    .INIT(32'h0133fecc))
    al_13048ea1 (
    .a(al_ebd95b94),
    .b(al_4690bf2e),
    .c(al_522428e2),
    .d(al_132ae268),
    .e(al_e8c5f626[4]),
    .o(al_7fea7bf));
  AL_MAP_LUT6 #(
    .EQN("(~B*(A*~(C)*D*~(E)*~(F)+~(A)*C*~(D)*E*~(F)+A*~(C)*D*E*~(F)+~(A)*C*D*E*~(F)+A*C*~(D)*~(E)*F+A*~(C)*D*~(E)*F+A*C*D*~(E)*F+~(A)*C*~(D)*E*F+A*C*~(D)*E*F+A*~(C)*D*E*F+~(A)*C*D*E*F+A*C*D*E*F))"),
    .INIT(64'h3230222012100200))
    al_aa3510f0 (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_d0555e9d[2]),
    .d(al_902efd00[15]),
    .e(al_902efd00[39]),
    .f(al_902efd00[47]),
    .o(al_f23520ad));
  AL_MAP_LUT5 #(
    .EQN("(~C*B*(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))"),
    .INIT(32'h0c080400))
    al_93d19f4b (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_d0555e9d[2]),
    .d(al_902efd00[23]),
    .e(al_902efd00[31]),
    .o(al_d48745aa));
  AL_MAP_LUT6 #(
    .EQN("(F*~(B*A*(C*~(D)*~(E)+~(C)*D*~(E)+C*D*~(E)+~(C)*~(D)*E+C*~(D)*E)))"),
    .INIT(64'hff77777f00000000))
    al_cba2ba8 (
    .a(al_7bce675b),
    .b(al_9e8909aa),
    .c(al_d0555e9d[0]),
    .d(al_d0555e9d[1]),
    .e(al_d0555e9d[2]),
    .f(al_902efd00[7]),
    .o(al_a8508f7c));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_8552c76c (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_902efd00[5]),
    .d(al_902efd00[13]),
    .e(al_902efd00[21]),
    .f(al_902efd00[29]),
    .o(al_29fafdbd));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_5c270cbf (
    .a(al_d0555e9d[0]),
    .b(al_902efd00[37]),
    .c(al_902efd00[45]),
    .o(al_a50e12e0));
  AL_MAP_LUT6 #(
    .EQN("~(A*~((~C*(E*~(F)*~(B)+E*F*~(B)+~(E)*F*B+E*F*B)))*~(D)+A*(~C*(E*~(F)*~(B)+E*F*~(B)+~(E)*F*B+E*F*B))*~(D)+~(A)*(~C*(E*~(F)*~(B)+E*F*~(B)+~(E)*F*B+E*F*B))*D+A*(~C*(E*~(F)*~(B)+E*F*~(B)+~(E)*F*B+E*F*B))*D)"),
    .INIT(64'hf055f355fc55ff55))
    al_df8ef082 (
    .a(al_2cc28140),
    .b(al_d0555e9d[0]),
    .c(al_d0555e9d[1]),
    .d(al_d0555e9d[2]),
    .e(al_902efd00[38]),
    .f(al_902efd00[46]),
    .o(al_f9f3df5f));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+~(A)*~(B)*~(C)*D*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+~(A)*B*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*D*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*C*D*E*~(F)+~(A)*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+~(A)*~(B)*C*D*~(E)*F+~(A)*B*C*D*~(E)*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F)"),
    .INIT(64'h00c05050ffcf5f5f))
    al_7575be31 (
    .a(al_29fafdbd),
    .b(al_a50e12e0),
    .c(al_132ae268),
    .d(al_d0555e9d[1]),
    .e(al_d0555e9d[2]),
    .f(al_902efd00[5]),
    .o(al_221dcd70));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_448661c6 (
    .a(al_d0555e9d[0]),
    .b(al_902efd00[34]),
    .c(al_902efd00[42]),
    .o(al_1af55219));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_7205fc52 (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_902efd00[2]),
    .d(al_902efd00[10]),
    .e(al_902efd00[18]),
    .f(al_902efd00[26]),
    .o(al_5e3e1251));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff3fafaf0030a0a0))
    al_27ca78dc (
    .a(al_5e3e1251),
    .b(al_1af55219),
    .c(al_132ae268),
    .d(al_d0555e9d[1]),
    .e(al_d0555e9d[2]),
    .f(al_902efd00[2]),
    .o(al_3a736cff[18]));
  AL_MAP_LUT6 #(
    .EQN("(~B*(A*~(C)*D*~(E)*~(F)+~(A)*C*~(D)*E*~(F)+A*~(C)*D*E*~(F)+~(A)*C*D*E*~(F)+A*C*~(D)*~(E)*F+A*~(C)*D*~(E)*F+A*C*D*~(E)*F+~(A)*C*~(D)*E*F+A*C*~(D)*E*F+A*~(C)*D*E*F+~(A)*C*D*E*F+A*C*D*E*F))"),
    .INIT(64'h3230222012100200))
    al_a8564136 (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_d0555e9d[2]),
    .d(al_902efd00[8]),
    .e(al_902efd00[32]),
    .f(al_902efd00[40]),
    .o(al_88de809d));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)*~(F)+A*~(B)*~(C)*~(D)*~(E)*~(F)+~(A)*B*~(C)*~(D)*~(E)*~(F)+A*B*~(C)*~(D)*~(E)*~(F)+~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*C*~(D)*~(E)*~(F)+~(A)*B*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*B*~(C)*D*~(E)*~(F)+A*B*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*~(B)*~(C)*~(D)*E*~(F)+A*~(B)*~(C)*~(D)*E*~(F)+A*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+A*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+~(A)*B*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F)"),
    .INIT(64'h32f336f73afb3eff))
    al_7ed116ad (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_d0555e9d[2]),
    .d(al_902efd00[0]),
    .e(al_902efd00[16]),
    .f(al_902efd00[24]),
    .o(al_d3c8ca1c));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_705ad0a9 (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_902efd00[3]),
    .d(al_902efd00[11]),
    .e(al_902efd00[19]),
    .f(al_902efd00[27]),
    .o(al_a51c3dde));
  AL_MAP_LUT6 #(
    .EQN("~(~A*~((~C*~(E*~(F)*~(B)+E*F*~(B)+~(E)*F*B+E*F*B)))*~(D)+~A*(~C*~(E*~(F)*~(B)+E*F*~(B)+~(E)*F*B+E*F*B))*~(D)+~(~A)*(~C*~(E*~(F)*~(B)+E*F*~(B)+~(E)*F*B+E*F*B))*D+~A*(~C*~(E*~(F)*~(B)+E*F*~(B)+~(E)*F*B+E*F*B))*D)"),
    .INIT(64'hffaafcaaf3aaf0aa))
    al_f27317b2 (
    .a(al_a51c3dde),
    .b(al_d0555e9d[0]),
    .c(al_d0555e9d[1]),
    .d(al_d0555e9d[2]),
    .e(al_902efd00[35]),
    .f(al_902efd00[43]),
    .o(al_c39b1824));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_8eb8b3a8 (
    .a(al_d0555e9d[0]),
    .b(al_902efd00[33]),
    .c(al_902efd00[41]),
    .o(al_b89e105d));
  AL_MAP_LUT6 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)*~(F)+A*~(B)*~(C)*D*~(E)*~(F)+~(A)*~(B)*C*D*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+~(A)*B*~(C)*~(D)*E*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+~(A)*B*C*~(D)*E*~(F)+A*~(B)*~(C)*D*E*~(F)+~(A)*B*~(C)*D*E*~(F)+~(A)*~(B)*C*D*E*~(F)+A*~(B)*C*D*E*~(F)+~(A)*B*C*D*E*~(F)+A*B*~(C)*~(D)*~(E)*F+~(A)*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+A*~(B)*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+~(A)*~(B)*C*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+~(A)*B*C*~(D)*E*F+A*B*C*~(D)*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hfedcba9876543210))
    al_bc7f0b1f (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_902efd00[1]),
    .d(al_902efd00[9]),
    .e(al_902efd00[17]),
    .f(al_902efd00[25]),
    .o(al_70936044));
  AL_MAP_LUT6 #(
    .EQN("(A*~(B)*C*~(D)*~(E)*~(F)+A*B*C*~(D)*~(E)*~(F)+A*~(B)*C*D*~(E)*~(F)+A*B*C*D*~(E)*~(F)+~(A)*~(B)*C*~(D)*E*~(F)+A*~(B)*C*~(D)*E*~(F)+~(A)*~(B)*~(C)*~(D)*~(E)*F+A*~(B)*~(C)*~(D)*~(E)*F+~(A)*B*~(C)*~(D)*~(E)*F+A*B*~(C)*~(D)*~(E)*F+A*~(B)*C*~(D)*~(E)*F+A*B*C*~(D)*~(E)*F+~(A)*~(B)*~(C)*D*~(E)*F+A*~(B)*~(C)*D*~(E)*F+~(A)*B*~(C)*D*~(E)*F+A*B*~(C)*D*~(E)*F+A*~(B)*C*D*~(E)*F+A*B*C*D*~(E)*F+~(A)*~(B)*~(C)*~(D)*E*F+A*~(B)*~(C)*~(D)*E*F+~(A)*B*~(C)*~(D)*E*F+A*B*~(C)*~(D)*E*F+~(A)*~(B)*C*~(D)*E*F+A*~(B)*C*~(D)*E*F+~(A)*~(B)*~(C)*D*E*F+A*~(B)*~(C)*D*E*F+~(A)*B*~(C)*D*E*F+A*B*~(C)*D*E*F+~(A)*~(B)*C*D*E*F+A*~(B)*C*D*E*F+~(A)*B*C*D*E*F+A*B*C*D*E*F)"),
    .INIT(64'hff3fafaf0030a0a0))
    al_b2829ef5 (
    .a(al_70936044),
    .b(al_b89e105d),
    .c(al_132ae268),
    .d(al_d0555e9d[1]),
    .e(al_d0555e9d[2]),
    .f(al_902efd00[1]),
    .o(al_3a736cff[17]));
  AL_MAP_LUT6 #(
    .EQN("(C@(~(A)*~(B)*~((E*D))*~(F)+A*~(B)*~((E*D))*~(F)+~(A)*B*~((E*D))*~(F)+~(A)*~(B)*(E*D)*~(F)+A*~(B)*(E*D)*~(F)+~(A)*B*(E*D)*~(F)+A*B*(E*D)*~(F)+~(A)*B*~((E*D))*F+~(A)*B*(E*D)*F))"),
    .INIT(64'hb4b4b4b40f878787))
    al_9481c889 (
    .a(al_c39b1824),
    .b(al_132ae268),
    .c(al_e8c5f626[3]),
    .d(al_d0555e9d[1]),
    .e(al_d0555e9d[2]),
    .f(al_902efd00[3]),
    .o(al_a2d9d6a));
  AL_MAP_LUT6 #(
    .EQN("(C@(~(A)*B*~((E*D))*~(F)+~(A)*B*(E*D)*~(F)+~(A)*~(B)*~((E*D))*F+A*~(B)*~((E*D))*F+~(A)*B*~((E*D))*F+~(A)*~(B)*(E*D)*F+A*~(B)*(E*D)*F+~(A)*B*(E*D)*F+A*B*(E*D)*F))"),
    .INIT(64'h0f878787b4b4b4b4))
    al_5bb97602 (
    .a(al_f9f3df5f),
    .b(al_132ae268),
    .c(al_e8c5f626[6]),
    .d(al_d0555e9d[1]),
    .e(al_d0555e9d[2]),
    .f(al_902efd00[6]),
    .o(al_ff09d078));
  AL_MAP_LUT5 #(
    .EQN("~(E@(~B*~(D*~(~C*~A))))"),
    .INIT(32'h0133fecc))
    al_d678aa25 (
    .a(al_f23520ad),
    .b(al_a8508f7c),
    .c(al_d48745aa),
    .d(al_132ae268),
    .e(al_e8c5f626[7]),
    .o(al_38f26a35));
  AL_MAP_LUT6 #(
    .EQN("(~B*~A*~(E@D)*~(F@C))"),
    .INIT(64'h1000001001000001))
    al_620b959f (
    .a(al_7fea7bf),
    .b(al_38f26a35),
    .c(al_3a736cff[18]),
    .d(al_3a736cff[17]),
    .e(al_e8c5f626[1]),
    .f(al_e8c5f626[2]),
    .o(al_a0e3e4ed));
  AL_MAP_LUT5 #(
    .EQN("(D@(~E*~((B*~A))*~(C)+~E*(B*~A)*~(C)+~(~E)*(B*~A)*C+~E*(B*~A)*C))"),
    .INIT(32'hbf40b04f))
    al_8fb034cf (
    .a(al_88de809d),
    .b(al_d3c8ca1c),
    .c(al_132ae268),
    .d(al_e8c5f626[0]),
    .e(al_902efd00[0]),
    .o(al_215b7b3d));
  AL_MAP_LUT3 #(
    .EQN("(C*(B@A))"),
    .INIT(8'h60))
    al_dbb48d8e (
    .a(al_221dcd70),
    .b(al_e8c5f626[5]),
    .c(al_d976dda9),
    .o(al_8d6efaba));
  AL_MAP_LUT6 #(
    .EQN("~(~F*~(E*D*C*~B*A))"),
    .INIT(64'hffffffff20000000))
    al_99e50bdf (
    .a(al_a0e3e4ed),
    .b(al_ff09d078),
    .c(al_a2d9d6a),
    .d(al_8d6efaba),
    .e(al_215b7b3d),
    .f(al_9b5719ae),
    .o(al_33c6f6));
  AL_MAP_LUT6 #(
    .EQN("(~B*(A*~(C)*D*~(E)*~(F)+~(A)*C*~(D)*E*~(F)+A*~(C)*D*E*~(F)+~(A)*C*D*E*~(F)+A*C*~(D)*~(E)*F+A*~(C)*D*~(E)*F+A*C*D*~(E)*F+~(A)*C*~(D)*E*F+A*C*~(D)*E*F+A*~(C)*D*E*F+~(A)*C*D*E*F+A*C*D*E*F))"),
    .INIT(64'h3230222012100200))
    al_4d1dd8ae (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_d0555e9d[2]),
    .d(al_902efd00[12]),
    .e(al_902efd00[36]),
    .f(al_902efd00[44]),
    .o(al_ebd95b94));
  AL_MAP_LUT5 #(
    .EQN("(~C*B*(D*~(E)*~(A)+D*E*~(A)+~(D)*E*A+D*E*A))"),
    .INIT(32'h0c080400))
    al_447a9367 (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_d0555e9d[2]),
    .d(al_902efd00[20]),
    .e(al_902efd00[28]),
    .o(al_522428e2));
  AL_MAP_LUT6 #(
    .EQN("(F*~(B*A*(C*~(D)*~(E)+~(C)*D*~(E)+C*D*~(E)+~(C)*~(D)*E+C*~(D)*E)))"),
    .INIT(64'hff77777f00000000))
    al_4a871a37 (
    .a(al_7bce675b),
    .b(al_9e8909aa),
    .c(al_d0555e9d[0]),
    .d(al_d0555e9d[1]),
    .e(al_d0555e9d[2]),
    .f(al_902efd00[4]),
    .o(al_4690bf2e));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_d091fda6 (
    .a(al_e8c5f626[1]),
    .b(al_e8c5f626[3]),
    .c(al_e8c5f626[5]),
    .o(al_68a14bd2));
  AL_MAP_LUT5 #(
    .EQN("(B*A*~(~D*~(~E*C)))"),
    .INIT(32'h88008880))
    al_59ce09d8 (
    .a(al_7bee3de4),
    .b(al_68a14bd2),
    .c(al_132ae268),
    .d(al_dbe2baa6),
    .e(al_30b5e311),
    .o(al_1c6db97d));
  AL_MAP_LUT6 #(
    .EQN("((E*~(D)*~((C*B))+E*D*~((C*B))+~(E)*D*(C*B)+E*D*(C*B))*~(~F*A))"),
    .INIT(64'hff3fc00055154000))
    al_e722f68b (
    .a(al_132ae268),
    .b(al_968fd17c),
    .c(al_d0555e9d[2]),
    .d(al_dbe2baa6),
    .e(al_7bec6b72),
    .f(al_30b5e311),
    .o(al_56997d45));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*C*B*~A)"),
    .INIT(64'h0000000000000040))
    al_a76da1ad (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_d0555e9d[2]),
    .d(al_dbe2baa6),
    .e(al_2110386e),
    .f(al_536b4576),
    .o(al_8e55a7af));
  AL_MAP_LUT6 #(
    .EQN("(~(B)*C*D*~(E)*~((~F*A))+~(B)*~(C)*~(D)*E*~((~F*A))+B*~(C)*~(D)*E*~((~F*A))+~(B)*C*~(D)*E*~((~F*A))+B*C*~(D)*E*~((~F*A))+~(B)*~(C)*D*E*~((~F*A))+B*~(C)*D*E*~((~F*A))+~(B)*C*D*E*~((~F*A))+B*C*D*E*~((~F*A))+~(B)*C*D*~(E)*(~F*A)+B*~(C)*~(D)*E*(~F*A)+~(B)*C*~(D)*E*(~F*A)+B*C*~(D)*E*(~F*A)+~(B)*~(C)*D*E*(~F*A)+B*~(C)*D*E*(~F*A)+~(B)*C*D*E*(~F*A)+B*C*D*E*(~F*A))"),
    .INIT(64'hffff3000fffd3000))
    al_1c093e97 (
    .a(al_132ae268),
    .b(al_d0555e9d[0]),
    .c(al_d0555e9d[1]),
    .d(al_d0555e9d[2]),
    .e(al_4596a396),
    .f(al_30b5e311),
    .o(al_9d9dbb20));
  AL_MAP_LUT6 #(
    .EQN("(A*~(~F*~E*~D*~C*B))"),
    .INIT(64'haaaaaaaaaaaaaaa2))
    al_4f7a09aa (
    .a(al_9d9dbb20),
    .b(al_8e55a7af),
    .c(al_8f15a934),
    .d(al_b5e36a9),
    .e(al_d976dda9),
    .f(al_3edda74b),
    .o(al_114295f1));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_188647e3 (
    .a(al_132ae268),
    .b(al_868a1cad[0]),
    .c(al_2408f449[8]),
    .o(al_40f6174[0]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_34108390 (
    .a(al_132ae268),
    .b(al_868a1cad[10]),
    .c(al_2408f449[18]),
    .o(al_40f6174[10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f0ba9b5 (
    .a(al_132ae268),
    .b(al_868a1cad[11]),
    .c(al_2408f449[19]),
    .o(al_40f6174[11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c4c4b2f2 (
    .a(al_132ae268),
    .b(al_868a1cad[12]),
    .c(al_2408f449[20]),
    .o(al_40f6174[12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_3a530990 (
    .a(al_132ae268),
    .b(al_868a1cad[13]),
    .c(al_2408f449[21]),
    .o(al_40f6174[13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_fc81f421 (
    .a(al_132ae268),
    .b(al_868a1cad[14]),
    .c(al_2408f449[22]),
    .o(al_40f6174[14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_7c5b49c5 (
    .a(al_132ae268),
    .b(al_868a1cad[15]),
    .c(al_2408f449[23]),
    .o(al_40f6174[15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e01428b6 (
    .a(al_132ae268),
    .b(al_868a1cad[16]),
    .c(al_2408f449[24]),
    .o(al_40f6174[16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1790332c (
    .a(al_132ae268),
    .b(al_868a1cad[17]),
    .c(al_2408f449[25]),
    .o(al_40f6174[17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_95987a97 (
    .a(al_132ae268),
    .b(al_868a1cad[18]),
    .c(al_2408f449[26]),
    .o(al_40f6174[18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d088cfd6 (
    .a(al_132ae268),
    .b(al_868a1cad[19]),
    .c(al_2408f449[27]),
    .o(al_40f6174[19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ec8e2d45 (
    .a(al_132ae268),
    .b(al_868a1cad[1]),
    .c(al_2408f449[9]),
    .o(al_40f6174[1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1fd9f289 (
    .a(al_132ae268),
    .b(al_868a1cad[20]),
    .c(al_2408f449[28]),
    .o(al_40f6174[20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8553b49b (
    .a(al_132ae268),
    .b(al_868a1cad[21]),
    .c(al_2408f449[29]),
    .o(al_40f6174[21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_6e38476a (
    .a(al_132ae268),
    .b(al_868a1cad[22]),
    .c(al_2408f449[30]),
    .o(al_40f6174[22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2f4d8714 (
    .a(al_132ae268),
    .b(al_868a1cad[23]),
    .c(al_2408f449[31]),
    .o(al_40f6174[23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b8cf30f4 (
    .a(al_132ae268),
    .b(al_868a1cad[24]),
    .c(al_2408f449[32]),
    .o(al_40f6174[24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_73cf2f5c (
    .a(al_132ae268),
    .b(al_868a1cad[25]),
    .c(al_2408f449[33]),
    .o(al_40f6174[25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9b307d1 (
    .a(al_132ae268),
    .b(al_868a1cad[26]),
    .c(al_2408f449[34]),
    .o(al_40f6174[26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8d6a1029 (
    .a(al_132ae268),
    .b(al_868a1cad[27]),
    .c(al_2408f449[35]),
    .o(al_40f6174[27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_da56d36d (
    .a(al_132ae268),
    .b(al_868a1cad[28]),
    .c(al_2408f449[36]),
    .o(al_40f6174[28]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d6dbaf55 (
    .a(al_132ae268),
    .b(al_868a1cad[29]),
    .c(al_2408f449[37]),
    .o(al_40f6174[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_90334166 (
    .a(al_132ae268),
    .b(al_868a1cad[2]),
    .c(al_2408f449[10]),
    .o(al_40f6174[2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_43f1371a (
    .a(al_132ae268),
    .b(al_868a1cad[30]),
    .c(al_2408f449[38]),
    .o(al_40f6174[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_881a9043 (
    .a(al_132ae268),
    .b(al_868a1cad[31]),
    .c(al_2408f449[39]),
    .o(al_40f6174[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b025e461 (
    .a(al_132ae268),
    .b(al_cd0aa0ee[0]),
    .c(al_2408f449[40]),
    .o(al_40f6174[32]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8771c034 (
    .a(al_132ae268),
    .b(al_cd0aa0ee[1]),
    .c(al_2408f449[41]),
    .o(al_40f6174[33]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f1c6c3b9 (
    .a(al_132ae268),
    .b(al_cd0aa0ee[2]),
    .c(al_2408f449[42]),
    .o(al_40f6174[34]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_5cc3e34b (
    .a(al_132ae268),
    .b(al_cd0aa0ee[3]),
    .c(al_2408f449[43]),
    .o(al_40f6174[35]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_25f391ce (
    .a(al_132ae268),
    .b(al_cd0aa0ee[4]),
    .c(al_2408f449[44]),
    .o(al_40f6174[36]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ca674493 (
    .a(al_132ae268),
    .b(al_cd0aa0ee[5]),
    .c(al_2408f449[45]),
    .o(al_40f6174[37]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e74b5503 (
    .a(al_132ae268),
    .b(al_cd0aa0ee[6]),
    .c(al_2408f449[46]),
    .o(al_40f6174[38]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_143371a (
    .a(al_132ae268),
    .b(al_cd0aa0ee[7]),
    .c(al_2408f449[47]),
    .o(al_40f6174[39]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_4c78ea1f (
    .a(al_132ae268),
    .b(al_868a1cad[3]),
    .c(al_2408f449[11]),
    .o(al_40f6174[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_815e71ca (
    .a(al_132ae268),
    .b(al_cd0aa0ee[8]),
    .o(al_40f6174[40]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_78d36b7b (
    .a(al_132ae268),
    .b(al_cd0aa0ee[9]),
    .o(al_40f6174[41]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_b0595909 (
    .a(al_132ae268),
    .b(al_cd0aa0ee[10]),
    .o(al_40f6174[42]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_3e96a041 (
    .a(al_132ae268),
    .b(al_cd0aa0ee[11]),
    .o(al_40f6174[43]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_69f87aea (
    .a(al_132ae268),
    .b(al_cd0aa0ee[12]),
    .o(al_40f6174[44]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_2e6cc269 (
    .a(al_132ae268),
    .b(al_cd0aa0ee[13]),
    .o(al_40f6174[45]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_b6d1f499 (
    .a(al_132ae268),
    .b(al_cd0aa0ee[14]),
    .o(al_40f6174[46]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_e945ae5c (
    .a(al_132ae268),
    .b(al_cd0aa0ee[15]),
    .o(al_40f6174[47]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a3f4d99a (
    .a(al_132ae268),
    .b(al_868a1cad[4]),
    .c(al_2408f449[12]),
    .o(al_40f6174[4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_60077b46 (
    .a(al_132ae268),
    .b(al_868a1cad[5]),
    .c(al_2408f449[13]),
    .o(al_40f6174[5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_5dcceb2f (
    .a(al_132ae268),
    .b(al_868a1cad[6]),
    .c(al_2408f449[14]),
    .o(al_40f6174[6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_7b3f2b12 (
    .a(al_132ae268),
    .b(al_868a1cad[7]),
    .c(al_2408f449[15]),
    .o(al_40f6174[7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9d9b1271 (
    .a(al_132ae268),
    .b(al_868a1cad[8]),
    .c(al_2408f449[16]),
    .o(al_40f6174[8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_225ed78c (
    .a(al_132ae268),
    .b(al_868a1cad[9]),
    .c(al_2408f449[17]),
    .o(al_40f6174[9]));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    al_9475c7cf (
    .a(al_e8c5f626[0]),
    .b(al_e8c5f626[7]),
    .c(al_2408f449[0]),
    .d(al_2408f449[7]),
    .o(al_f16b3d6d));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    al_a0cb837f (
    .a(al_f16b3d6d),
    .b(al_e8c5f626[3]),
    .c(al_e8c5f626[5]),
    .d(al_2408f449[3]),
    .e(al_2408f449[5]),
    .o(al_49c7fc0e));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    al_bb903191 (
    .a(al_e8c5f626[2]),
    .b(al_e8c5f626[4]),
    .c(al_2408f449[2]),
    .d(al_2408f449[4]),
    .o(al_113d1401));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    al_a0de75ee (
    .a(al_113d1401),
    .b(al_e8c5f626[1]),
    .c(al_e8c5f626[6]),
    .d(al_2408f449[1]),
    .e(al_2408f449[6]),
    .o(al_8e145e50));
  AL_MAP_LUT5 #(
    .EQN("(B*A*~(~D*~(~E*C)))"),
    .INIT(32'h88008880))
    al_5e86ff7c (
    .a(al_49c7fc0e),
    .b(al_8e145e50),
    .c(al_132ae268),
    .d(al_2110386e),
    .e(al_30b5e311),
    .o(al_982b355d));
  AL_MAP_LUT6 #(
    .EQN("((E*~(D)*~((C*B))+E*D*~((C*B))+~(E)*D*(C*B)+E*D*(C*B))*~(~F*A))"),
    .INIT(64'hff3fc00055154000))
    al_46f88da0 (
    .a(al_132ae268),
    .b(al_968fd17c),
    .c(al_d0555e9d[2]),
    .d(al_2110386e),
    .e(al_88c53423),
    .f(al_30b5e311),
    .o(al_4efdb29f));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_a10ebaec (
    .a(al_132ae268),
    .b(al_2bdcc449[8]),
    .c(al_49a90ce2[0]),
    .o(al_f0cac652[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_eb07cf02 (
    .a(al_132ae268),
    .b(al_2bdcc449[18]),
    .c(al_49a90ce2[10]),
    .o(al_f0cac652[10]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_d8df1e13 (
    .a(al_132ae268),
    .b(al_2bdcc449[19]),
    .c(al_49a90ce2[11]),
    .o(al_f0cac652[11]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_3ca5e072 (
    .a(al_132ae268),
    .b(al_2bdcc449[20]),
    .c(al_49a90ce2[12]),
    .o(al_f0cac652[12]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_c303f104 (
    .a(al_132ae268),
    .b(al_2bdcc449[21]),
    .c(al_49a90ce2[13]),
    .o(al_f0cac652[13]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_c5d6fe17 (
    .a(al_132ae268),
    .b(al_2bdcc449[22]),
    .c(al_49a90ce2[14]),
    .o(al_f0cac652[14]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_683e81a3 (
    .a(al_132ae268),
    .b(al_2bdcc449[23]),
    .c(al_49a90ce2[15]),
    .o(al_f0cac652[15]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_fcf481b0 (
    .a(al_132ae268),
    .b(al_2bdcc449[24]),
    .c(al_49a90ce2[16]),
    .o(al_f0cac652[16]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_fa960790 (
    .a(al_132ae268),
    .b(al_2bdcc449[25]),
    .c(al_49a90ce2[17]),
    .o(al_f0cac652[17]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_a7db0aef (
    .a(al_132ae268),
    .b(al_2bdcc449[26]),
    .c(al_49a90ce2[18]),
    .o(al_f0cac652[18]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_d8d9afdd (
    .a(al_132ae268),
    .b(al_2bdcc449[27]),
    .c(al_49a90ce2[19]),
    .o(al_f0cac652[19]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_c51cd03f (
    .a(al_132ae268),
    .b(al_2bdcc449[9]),
    .c(al_49a90ce2[1]),
    .o(al_f0cac652[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_c2484409 (
    .a(al_132ae268),
    .b(al_2bdcc449[28]),
    .c(al_49a90ce2[20]),
    .o(al_f0cac652[20]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_38f91704 (
    .a(al_132ae268),
    .b(al_2bdcc449[29]),
    .c(al_49a90ce2[21]),
    .o(al_f0cac652[21]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_3c3e34c7 (
    .a(al_132ae268),
    .b(al_2bdcc449[30]),
    .c(al_49a90ce2[22]),
    .o(al_f0cac652[22]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_377335df (
    .a(al_132ae268),
    .b(al_2bdcc449[31]),
    .c(al_49a90ce2[23]),
    .o(al_f0cac652[23]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_4a4a487d (
    .a(al_132ae268),
    .b(al_2bdcc449[32]),
    .c(al_49a90ce2[24]),
    .o(al_f0cac652[24]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_f4500095 (
    .a(al_132ae268),
    .b(al_2bdcc449[33]),
    .c(al_49a90ce2[25]),
    .o(al_f0cac652[25]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_f2eb511e (
    .a(al_132ae268),
    .b(al_2bdcc449[34]),
    .c(al_49a90ce2[26]),
    .o(al_f0cac652[26]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_2607991e (
    .a(al_132ae268),
    .b(al_2bdcc449[35]),
    .c(al_49a90ce2[27]),
    .o(al_f0cac652[27]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_810512dd (
    .a(al_132ae268),
    .b(al_2bdcc449[36]),
    .c(al_49a90ce2[28]),
    .o(al_f0cac652[28]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_358991b (
    .a(al_132ae268),
    .b(al_2bdcc449[37]),
    .c(al_49a90ce2[29]),
    .o(al_f0cac652[29]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_2e03fcd3 (
    .a(al_132ae268),
    .b(al_2bdcc449[10]),
    .c(al_49a90ce2[2]),
    .o(al_f0cac652[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_dc297c23 (
    .a(al_132ae268),
    .b(al_2bdcc449[38]),
    .c(al_49a90ce2[30]),
    .o(al_f0cac652[30]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_62b0bcdc (
    .a(al_132ae268),
    .b(al_2bdcc449[39]),
    .c(al_49a90ce2[31]),
    .o(al_f0cac652[31]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_96cb37b8 (
    .a(al_132ae268),
    .b(al_2bdcc449[40]),
    .c(al_49a90ce2[32]),
    .o(al_f0cac652[32]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_decb0334 (
    .a(al_132ae268),
    .b(al_2bdcc449[41]),
    .c(al_49a90ce2[33]),
    .o(al_f0cac652[33]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_9b42e552 (
    .a(al_132ae268),
    .b(al_2bdcc449[42]),
    .c(al_49a90ce2[34]),
    .o(al_f0cac652[34]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_9f32d1ee (
    .a(al_132ae268),
    .b(al_2bdcc449[43]),
    .c(al_49a90ce2[35]),
    .o(al_f0cac652[35]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_55353a59 (
    .a(al_132ae268),
    .b(al_2bdcc449[44]),
    .c(al_49a90ce2[36]),
    .o(al_f0cac652[36]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_639fbaa1 (
    .a(al_132ae268),
    .b(al_2bdcc449[45]),
    .c(al_49a90ce2[37]),
    .o(al_f0cac652[37]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_6e6768b5 (
    .a(al_132ae268),
    .b(al_2bdcc449[46]),
    .c(al_49a90ce2[38]),
    .o(al_f0cac652[38]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_e00fa476 (
    .a(al_132ae268),
    .b(al_2bdcc449[47]),
    .c(al_49a90ce2[39]),
    .o(al_f0cac652[39]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_61947c9a (
    .a(al_132ae268),
    .b(al_2bdcc449[11]),
    .c(al_49a90ce2[3]),
    .o(al_f0cac652[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_ccb9481f (
    .a(al_132ae268),
    .b(al_49a90ce2[40]),
    .o(al_f0cac652[40]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_db7f9207 (
    .a(al_132ae268),
    .b(al_49a90ce2[41]),
    .o(al_f0cac652[41]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_4f3dfeb3 (
    .a(al_132ae268),
    .b(al_49a90ce2[42]),
    .o(al_f0cac652[42]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_dfde759b (
    .a(al_132ae268),
    .b(al_49a90ce2[43]),
    .o(al_f0cac652[43]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_cff3a8bb (
    .a(al_132ae268),
    .b(al_49a90ce2[44]),
    .o(al_f0cac652[44]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_c4270e05 (
    .a(al_132ae268),
    .b(al_49a90ce2[45]),
    .o(al_f0cac652[45]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_4a2021c1 (
    .a(al_132ae268),
    .b(al_49a90ce2[46]),
    .o(al_f0cac652[46]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_6fa38b7a (
    .a(al_132ae268),
    .b(al_49a90ce2[47]),
    .o(al_f0cac652[47]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_ecbd335f (
    .a(al_132ae268),
    .b(al_2bdcc449[12]),
    .c(al_49a90ce2[4]),
    .o(al_f0cac652[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_9a3cb4ea (
    .a(al_132ae268),
    .b(al_2bdcc449[13]),
    .c(al_49a90ce2[5]),
    .o(al_f0cac652[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_ccee842b (
    .a(al_132ae268),
    .b(al_2bdcc449[14]),
    .c(al_49a90ce2[6]),
    .o(al_f0cac652[6]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_ace9f52 (
    .a(al_132ae268),
    .b(al_2bdcc449[15]),
    .c(al_49a90ce2[7]),
    .o(al_f0cac652[7]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_4485624e (
    .a(al_132ae268),
    .b(al_2bdcc449[16]),
    .c(al_49a90ce2[8]),
    .o(al_f0cac652[8]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_ac1e6add (
    .a(al_132ae268),
    .b(al_2bdcc449[17]),
    .c(al_49a90ce2[9]),
    .o(al_f0cac652[9]));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    al_8c300dd6 (
    .a(al_e8c5f626[2]),
    .b(al_e8c5f626[7]),
    .c(al_2bdcc449[2]),
    .d(al_2bdcc449[7]),
    .o(al_56b3d928));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    al_5510d5c5 (
    .a(al_56b3d928),
    .b(al_e8c5f626[4]),
    .c(al_e8c5f626[5]),
    .d(al_2bdcc449[4]),
    .e(al_2bdcc449[5]),
    .o(al_66d47dbf));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    al_d55b72d0 (
    .a(al_e8c5f626[0]),
    .b(al_e8c5f626[1]),
    .c(al_2bdcc449[0]),
    .d(al_2bdcc449[1]),
    .o(al_dc21b291));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    al_db1dc4a6 (
    .a(al_dc21b291),
    .b(al_e8c5f626[3]),
    .c(al_e8c5f626[6]),
    .d(al_2bdcc449[3]),
    .e(al_2bdcc449[6]),
    .o(al_db67c2f5));
  AL_MAP_LUT5 #(
    .EQN("(B*A*~(~D*~(~E*C)))"),
    .INIT(32'h88008880))
    al_bcba5d98 (
    .a(al_66d47dbf),
    .b(al_db67c2f5),
    .c(al_132ae268),
    .d(al_536b4576),
    .e(al_30b5e311),
    .o(al_3e178366));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    al_798b6f6c (
    .a(al_82716c38[4]),
    .b(al_82716c38[5]),
    .c(al_82716c38[6]),
    .d(al_82716c38[7]),
    .o(al_e4f9c44c));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_b451064 (
    .a(al_d23bd93a),
    .b(s_axi_wdata[0]),
    .c(unicast_addr[0]),
    .d(al_81344cef),
    .e(al_49a90ce2[0]),
    .o(al_9db0b0fa[0]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_8921eae1 (
    .a(al_d23bd93a),
    .b(s_axi_wdata[10]),
    .c(unicast_addr[10]),
    .d(al_81344cef),
    .e(al_49a90ce2[10]),
    .o(al_9db0b0fa[10]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_124ab9ab (
    .a(al_d23bd93a),
    .b(s_axi_wdata[11]),
    .c(unicast_addr[11]),
    .d(al_81344cef),
    .e(al_49a90ce2[11]),
    .o(al_9db0b0fa[11]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_ba384718 (
    .a(al_d23bd93a),
    .b(s_axi_wdata[12]),
    .c(unicast_addr[12]),
    .d(al_81344cef),
    .e(al_49a90ce2[12]),
    .o(al_9db0b0fa[12]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_44ef27a6 (
    .a(al_d23bd93a),
    .b(s_axi_wdata[13]),
    .c(unicast_addr[13]),
    .d(al_81344cef),
    .e(al_49a90ce2[13]),
    .o(al_9db0b0fa[13]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_b75ed0b8 (
    .a(al_d23bd93a),
    .b(s_axi_wdata[14]),
    .c(unicast_addr[14]),
    .d(al_81344cef),
    .e(al_49a90ce2[14]),
    .o(al_9db0b0fa[14]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_f14e7b71 (
    .a(al_d23bd93a),
    .b(s_axi_wdata[15]),
    .c(unicast_addr[15]),
    .d(al_81344cef),
    .e(al_49a90ce2[15]),
    .o(al_9db0b0fa[15]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_92e952c2 (
    .a(al_d23bd93a),
    .b(s_axi_wdata[16]),
    .c(unicast_addr[16]),
    .d(al_81344cef),
    .e(al_49a90ce2[16]),
    .o(al_9db0b0fa[16]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_f01ba3d2 (
    .a(al_d23bd93a),
    .b(s_axi_wdata[17]),
    .c(unicast_addr[17]),
    .d(al_81344cef),
    .e(al_49a90ce2[17]),
    .o(al_9db0b0fa[17]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_d5a83ec8 (
    .a(al_d23bd93a),
    .b(s_axi_wdata[18]),
    .c(unicast_addr[18]),
    .d(al_81344cef),
    .e(al_49a90ce2[18]),
    .o(al_9db0b0fa[18]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_d83269ae (
    .a(al_d23bd93a),
    .b(s_axi_wdata[19]),
    .c(unicast_addr[19]),
    .d(al_81344cef),
    .e(al_49a90ce2[19]),
    .o(al_9db0b0fa[19]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_34a77175 (
    .a(al_d23bd93a),
    .b(s_axi_wdata[1]),
    .c(unicast_addr[1]),
    .d(al_81344cef),
    .e(al_49a90ce2[1]),
    .o(al_9db0b0fa[1]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_246ca3a6 (
    .a(al_d23bd93a),
    .b(s_axi_wdata[20]),
    .c(unicast_addr[20]),
    .d(al_81344cef),
    .e(al_49a90ce2[20]),
    .o(al_9db0b0fa[20]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_8392aced (
    .a(al_d23bd93a),
    .b(s_axi_wdata[21]),
    .c(unicast_addr[21]),
    .d(al_81344cef),
    .e(al_49a90ce2[21]),
    .o(al_9db0b0fa[21]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_3cc9c657 (
    .a(al_d23bd93a),
    .b(s_axi_wdata[22]),
    .c(unicast_addr[22]),
    .d(al_81344cef),
    .e(al_49a90ce2[22]),
    .o(al_9db0b0fa[22]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_889ae054 (
    .a(al_d23bd93a),
    .b(s_axi_wdata[23]),
    .c(unicast_addr[23]),
    .d(al_81344cef),
    .e(al_49a90ce2[23]),
    .o(al_9db0b0fa[23]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_8b822842 (
    .a(al_d23bd93a),
    .b(s_axi_wdata[24]),
    .c(unicast_addr[24]),
    .d(al_81344cef),
    .e(al_49a90ce2[24]),
    .o(al_9db0b0fa[24]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_9d6b5c2b (
    .a(al_d23bd93a),
    .b(s_axi_wdata[25]),
    .c(unicast_addr[25]),
    .d(al_81344cef),
    .e(al_49a90ce2[25]),
    .o(al_9db0b0fa[25]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_f6d0b11c (
    .a(al_d23bd93a),
    .b(s_axi_wdata[26]),
    .c(unicast_addr[26]),
    .d(al_81344cef),
    .e(al_49a90ce2[26]),
    .o(al_9db0b0fa[26]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_5a83f853 (
    .a(al_d23bd93a),
    .b(s_axi_wdata[27]),
    .c(unicast_addr[27]),
    .d(al_81344cef),
    .e(al_49a90ce2[27]),
    .o(al_9db0b0fa[27]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_3d69c270 (
    .a(al_d23bd93a),
    .b(s_axi_wdata[28]),
    .c(unicast_addr[28]),
    .d(al_81344cef),
    .e(al_49a90ce2[28]),
    .o(al_9db0b0fa[28]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_e83960ce (
    .a(al_d23bd93a),
    .b(s_axi_wdata[29]),
    .c(unicast_addr[29]),
    .d(al_81344cef),
    .e(al_49a90ce2[29]),
    .o(al_9db0b0fa[29]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_a0d4091b (
    .a(al_d23bd93a),
    .b(s_axi_wdata[2]),
    .c(unicast_addr[2]),
    .d(al_81344cef),
    .e(al_49a90ce2[2]),
    .o(al_9db0b0fa[2]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    al_4a68f543 (
    .a(al_5df5c44f),
    .b(al_13660933[0]),
    .c(al_13660933[1]),
    .d(al_13660933[2]),
    .e(al_13660933[3]),
    .o(al_cf696ef0));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_c6a0ff5e (
    .a(al_cf696ef0),
    .b(al_41ffdcd4),
    .c(al_13660933[4]),
    .d(al_13660933[5]),
    .o(al_d23bd93a));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_f3b11212 (
    .a(al_d23bd93a),
    .b(s_axi_wdata[30]),
    .c(unicast_addr[30]),
    .d(al_81344cef),
    .e(al_49a90ce2[30]),
    .o(al_9db0b0fa[30]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_bda9f2e0 (
    .a(al_d23bd93a),
    .b(s_axi_wdata[31]),
    .c(unicast_addr[31]),
    .d(al_81344cef),
    .e(al_49a90ce2[31]),
    .o(al_9db0b0fa[31]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_1d015712 (
    .a(al_f7638b94),
    .b(s_axi_wdata[0]),
    .c(unicast_addr[32]),
    .d(al_81344cef),
    .e(al_49a90ce2[32]),
    .o(al_9db0b0fa[32]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_b7a10340 (
    .a(al_f7638b94),
    .b(s_axi_wdata[1]),
    .c(unicast_addr[33]),
    .d(al_81344cef),
    .e(al_49a90ce2[33]),
    .o(al_9db0b0fa[33]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_3fd51d3b (
    .a(al_f7638b94),
    .b(s_axi_wdata[2]),
    .c(unicast_addr[34]),
    .d(al_81344cef),
    .e(al_49a90ce2[34]),
    .o(al_9db0b0fa[34]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_56043e0c (
    .a(al_f7638b94),
    .b(s_axi_wdata[3]),
    .c(unicast_addr[35]),
    .d(al_81344cef),
    .e(al_49a90ce2[35]),
    .o(al_9db0b0fa[35]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_c435b48e (
    .a(al_f7638b94),
    .b(s_axi_wdata[4]),
    .c(unicast_addr[36]),
    .d(al_81344cef),
    .e(al_49a90ce2[36]),
    .o(al_9db0b0fa[36]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_b76181bc (
    .a(al_f7638b94),
    .b(s_axi_wdata[5]),
    .c(unicast_addr[37]),
    .d(al_81344cef),
    .e(al_49a90ce2[37]),
    .o(al_9db0b0fa[37]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_89fc5163 (
    .a(al_f7638b94),
    .b(s_axi_wdata[6]),
    .c(unicast_addr[38]),
    .d(al_81344cef),
    .e(al_49a90ce2[38]),
    .o(al_9db0b0fa[38]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_fa7ce057 (
    .a(al_f7638b94),
    .b(s_axi_wdata[7]),
    .c(unicast_addr[39]),
    .d(al_81344cef),
    .e(al_49a90ce2[39]),
    .o(al_9db0b0fa[39]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_785996d5 (
    .a(al_d23bd93a),
    .b(s_axi_wdata[3]),
    .c(unicast_addr[3]),
    .d(al_81344cef),
    .e(al_49a90ce2[3]),
    .o(al_9db0b0fa[3]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_1260e293 (
    .a(al_f7638b94),
    .b(s_axi_wdata[8]),
    .c(unicast_addr[40]),
    .d(al_81344cef),
    .e(al_49a90ce2[40]),
    .o(al_9db0b0fa[40]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_56c7736f (
    .a(al_f7638b94),
    .b(s_axi_wdata[9]),
    .c(unicast_addr[41]),
    .d(al_81344cef),
    .e(al_49a90ce2[41]),
    .o(al_9db0b0fa[41]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_4c92f5de (
    .a(al_f7638b94),
    .b(s_axi_wdata[10]),
    .c(unicast_addr[42]),
    .d(al_81344cef),
    .e(al_49a90ce2[42]),
    .o(al_9db0b0fa[42]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_5c3b6bcd (
    .a(al_f7638b94),
    .b(s_axi_wdata[11]),
    .c(unicast_addr[43]),
    .d(al_81344cef),
    .e(al_49a90ce2[43]),
    .o(al_9db0b0fa[43]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_59939512 (
    .a(al_f7638b94),
    .b(s_axi_wdata[12]),
    .c(unicast_addr[44]),
    .d(al_81344cef),
    .e(al_49a90ce2[44]),
    .o(al_9db0b0fa[44]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_8b167973 (
    .a(al_f7638b94),
    .b(s_axi_wdata[13]),
    .c(unicast_addr[45]),
    .d(al_81344cef),
    .e(al_49a90ce2[45]),
    .o(al_9db0b0fa[45]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_e7cea1fd (
    .a(al_7afe69f4),
    .b(al_5df5c44f),
    .c(al_13660933[2]),
    .d(al_13660933[3]),
    .o(al_f7638b94));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_39acbb54 (
    .a(al_f7638b94),
    .b(s_axi_wdata[14]),
    .c(unicast_addr[46]),
    .d(al_81344cef),
    .e(al_49a90ce2[46]),
    .o(al_9db0b0fa[46]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_276f1208 (
    .a(al_f7638b94),
    .b(s_axi_wdata[15]),
    .c(unicast_addr[47]),
    .d(al_81344cef),
    .e(al_49a90ce2[47]),
    .o(al_9db0b0fa[47]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_9b2549e4 (
    .a(al_d23bd93a),
    .b(s_axi_wdata[4]),
    .c(unicast_addr[4]),
    .d(al_81344cef),
    .e(al_49a90ce2[4]),
    .o(al_9db0b0fa[4]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_d0d51cbb (
    .a(al_d23bd93a),
    .b(s_axi_wdata[5]),
    .c(unicast_addr[5]),
    .d(al_81344cef),
    .e(al_49a90ce2[5]),
    .o(al_9db0b0fa[5]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_cd9ca72c (
    .a(al_d23bd93a),
    .b(s_axi_wdata[6]),
    .c(unicast_addr[6]),
    .d(al_81344cef),
    .e(al_49a90ce2[6]),
    .o(al_9db0b0fa[6]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_38b4d90f (
    .a(al_d23bd93a),
    .b(s_axi_wdata[7]),
    .c(unicast_addr[7]),
    .d(al_81344cef),
    .e(al_49a90ce2[7]),
    .o(al_9db0b0fa[7]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_66c31acd (
    .a(al_d23bd93a),
    .b(s_axi_wdata[8]),
    .c(unicast_addr[8]),
    .d(al_81344cef),
    .e(al_49a90ce2[8]),
    .o(al_9db0b0fa[8]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*~(C)*~(D)+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*~(D)+~((E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))*C*D+(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A)*C*D)"),
    .INIT(32'hf0ddf088))
    al_58af0c2d (
    .a(al_d23bd93a),
    .b(s_axi_wdata[9]),
    .c(unicast_addr[9]),
    .d(al_81344cef),
    .e(al_49a90ce2[9]),
    .o(al_9db0b0fa[9]));
  AL_MAP_LUT5 #(
    .EQN("(A*~((~(~D*~C)*~B))*~(E)+~(A)*(~(~D*~C)*~B)*~(E)+A*(~(~D*~C)*~B)*~(E)+A*(~(~D*~C)*~B)*E)"),
    .INIT(32'h2220bbba))
    al_7c232414 (
    .a(al_132ae268),
    .b(al_d0555e9d[0]),
    .c(al_d0555e9d[1]),
    .d(al_d0555e9d[2]),
    .e(al_30b5e311),
    .o(al_7e8a07be[0]));
  AL_MAP_LUT4 #(
    .EQN("((C@B)*~(D@A))"),
    .INIT(16'h2814))
    al_c3e2ffaa (
    .a(al_132ae268),
    .b(al_d0555e9d[0]),
    .c(al_d0555e9d[1]),
    .d(al_30b5e311),
    .o(al_7e8a07be[1]));
  AL_MAP_LUT5 #(
    .EQN("((D@(C*B))*~(E@A))"),
    .INIT(32'h2a801540))
    al_ff81820b (
    .a(al_132ae268),
    .b(al_d0555e9d[0]),
    .c(al_d0555e9d[1]),
    .d(al_d0555e9d[2]),
    .e(al_30b5e311),
    .o(al_7e8a07be[2]));
  AL_DFF_X al_42545c79 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_982b355d),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_2110386e));
  AL_DFF_X al_d00dfd58 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_4efdb29f),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_88c53423));
  AL_DFF_X al_c953fa3d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_62d97d99),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad22e376));
  AL_MAP_LUT5 #(
    .EQN("(~C*(E*~(D)*~((B*A))+E*D*~((B*A))+~(E)*D*(B*A)+E*D*(B*A)))"),
    .INIT(32'h0f070800))
    al_c1dd2b0f (
    .a(al_473186ca),
    .b(rx_clk_en),
    .c(al_ff9a7266),
    .d(al_a9406400),
    .e(al_ad22e376),
    .o(al_62d97d99));
  AL_DFF_X al_85a91f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_7e8a07be[0]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_d0555e9d[0]));
  AL_DFF_X al_cad329bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_7e8a07be[1]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_d0555e9d[1]));
  AL_DFF_X al_ce44cbb6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_7e8a07be[2]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_d0555e9d[2]));
  AL_DFF_X al_edfcc04c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[0]),
    .en(al_8f82c712),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[0]));
  AL_DFF_X al_24345f6f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[9]),
    .en(al_8f82c712),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[9]));
  AL_DFF_X al_28cd96e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[10]),
    .en(al_8f82c712),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[10]));
  AL_DFF_X al_22cfaf24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[11]),
    .en(al_8f82c712),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[11]));
  AL_DFF_X al_19d967c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[12]),
    .en(al_8f82c712),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[12]));
  AL_DFF_X al_5b71aff3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[13]),
    .en(al_8f82c712),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[13]));
  AL_DFF_X al_5fc792a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[14]),
    .en(al_8f82c712),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[14]));
  AL_DFF_X al_cecf5c1b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[15]),
    .en(al_8f82c712),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[15]));
  AL_DFF_X al_2fc73c6d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[16]),
    .en(al_8f82c712),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[16]));
  AL_DFF_X al_65d0a199 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[17]),
    .en(al_8f82c712),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[17]));
  AL_DFF_X al_14eef1ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[18]),
    .en(al_8f82c712),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[18]));
  AL_DFF_X al_d6ff79c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[1]),
    .en(al_8f82c712),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[1]));
  AL_DFF_X al_e47d66e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[19]),
    .en(al_8f82c712),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[19]));
  AL_DFF_X al_43acd35f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[20]),
    .en(al_8f82c712),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[20]));
  AL_DFF_X al_de250307 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[21]),
    .en(al_8f82c712),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[21]));
  AL_DFF_X al_32a52838 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[22]),
    .en(al_8f82c712),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[22]));
  AL_DFF_X al_8fe85d65 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[23]),
    .en(al_8f82c712),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[23]));
  AL_DFF_X al_ec1b4a4d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[24]),
    .en(al_8f82c712),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[24]));
  AL_DFF_X al_ecd47d6c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[25]),
    .en(al_8f82c712),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[25]));
  AL_DFF_X al_25c8f101 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[26]),
    .en(al_8f82c712),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[26]));
  AL_DFF_X al_cf7cd1a1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[27]),
    .en(al_8f82c712),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[27]));
  AL_DFF_X al_c2042f4d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[28]),
    .en(al_8f82c712),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[28]));
  AL_DFF_X al_5d043718 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[2]),
    .en(al_8f82c712),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[2]));
  AL_DFF_X al_18aa9b96 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[29]),
    .en(al_8f82c712),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[29]));
  AL_DFF_X al_cea465cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[30]),
    .en(al_8f82c712),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[30]));
  AL_DFF_X al_90c7c05f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[31]),
    .en(al_8f82c712),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[31]));
  AL_DFF_X al_2df377fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[0]),
    .en(al_71f17e1a),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[32]));
  AL_DFF_X al_b792488e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[1]),
    .en(al_71f17e1a),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[33]));
  AL_DFF_X al_2d677933 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[2]),
    .en(al_71f17e1a),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[34]));
  AL_DFF_X al_70f52f4e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[3]),
    .en(al_71f17e1a),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[35]));
  AL_DFF_X al_172ff953 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[4]),
    .en(al_71f17e1a),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[36]));
  AL_DFF_X al_2ffd93ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[5]),
    .en(al_71f17e1a),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[37]));
  AL_DFF_X al_2caf7fb7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[6]),
    .en(al_71f17e1a),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[38]));
  AL_DFF_X al_ec53ec7b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[3]),
    .en(al_8f82c712),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[3]));
  AL_DFF_X al_e7ca7957 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[7]),
    .en(al_71f17e1a),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[39]));
  AL_DFF_X al_be6d0b3c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[8]),
    .en(al_71f17e1a),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[40]));
  AL_DFF_X al_4a8b88d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[9]),
    .en(al_71f17e1a),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[41]));
  AL_DFF_X al_a43e4a54 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[10]),
    .en(al_71f17e1a),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[42]));
  AL_DFF_X al_de1e960b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[11]),
    .en(al_71f17e1a),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[43]));
  AL_DFF_X al_df7dc927 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[12]),
    .en(al_71f17e1a),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[44]));
  AL_DFF_X al_6af9af6f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[13]),
    .en(al_71f17e1a),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[45]));
  AL_DFF_X al_4280c84e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[14]),
    .en(al_71f17e1a),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[46]));
  AL_DFF_X al_a119eda6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[15]),
    .en(al_71f17e1a),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[47]));
  AL_DFF_X al_5832c5e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[16]),
    .en(al_71f17e1a),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[48]));
  AL_DFF_X al_3035e536 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[4]),
    .en(al_8f82c712),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[4]));
  AL_DFF_X al_303c54d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[17]),
    .en(al_71f17e1a),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[49]));
  AL_DFF_X al_fc3ebbb0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[18]),
    .en(al_71f17e1a),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[50]));
  AL_DFF_X al_c5476c96 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[19]),
    .en(al_71f17e1a),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[51]));
  AL_DFF_X al_4fa2e98b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[20]),
    .en(al_71f17e1a),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[52]));
  AL_DFF_X al_45b76947 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[21]),
    .en(al_71f17e1a),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[53]));
  AL_DFF_X al_d6bae0ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[22]),
    .en(al_71f17e1a),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[54]));
  AL_DFF_X al_3f369ec2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[23]),
    .en(al_71f17e1a),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[55]));
  AL_DFF_X al_b29c3483 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[24]),
    .en(al_71f17e1a),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[56]));
  AL_DFF_X al_24ca2aac (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[25]),
    .en(al_71f17e1a),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[57]));
  AL_DFF_X al_614df6af (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[26]),
    .en(al_71f17e1a),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[58]));
  AL_DFF_X al_20c389f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[5]),
    .en(al_8f82c712),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[5]));
  AL_DFF_X al_e4a1409e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[27]),
    .en(al_71f17e1a),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[59]));
  AL_DFF_X al_4bc283c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[28]),
    .en(al_71f17e1a),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[60]));
  AL_DFF_X al_5bb04a17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[29]),
    .en(al_71f17e1a),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[61]));
  AL_DFF_X al_c25655c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[30]),
    .en(al_71f17e1a),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[62]));
  AL_DFF_X al_3b2955bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[31]),
    .en(al_71f17e1a),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[63]));
  AL_DFF_X al_b30cbf5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[6]),
    .en(al_8f82c712),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[6]));
  AL_DFF_X al_4293aa44 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[7]),
    .en(al_8f82c712),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[7]));
  AL_DFF_X al_cce5ec27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[8]),
    .en(al_8f82c712),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_902efd00[8]));
  AL_DFF_X al_76ee72de (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[0]),
    .en(al_82faa065),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[0]));
  AL_DFF_X al_88b6b6ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[9]),
    .en(al_82faa065),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[9]));
  AL_DFF_X al_2679048f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[10]),
    .en(al_82faa065),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[10]));
  AL_DFF_X al_7852959f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[11]),
    .en(al_82faa065),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[11]));
  AL_DFF_X al_299a02e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[12]),
    .en(al_82faa065),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[12]));
  AL_DFF_X al_c0b5f642 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[13]),
    .en(al_82faa065),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[13]));
  AL_DFF_X al_4a1f4d14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[14]),
    .en(al_82faa065),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[14]));
  AL_DFF_X al_2437913b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[15]),
    .en(al_82faa065),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[15]));
  AL_DFF_X al_23bfdb97 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[16]),
    .en(al_82faa065),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[16]));
  AL_DFF_X al_fdc08dee (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[17]),
    .en(al_82faa065),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[17]));
  AL_DFF_X al_fcfa6d0e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[18]),
    .en(al_82faa065),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[18]));
  AL_DFF_X al_1d8665d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[1]),
    .en(al_82faa065),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[1]));
  AL_DFF_X al_93230eeb (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[19]),
    .en(al_82faa065),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[19]));
  AL_DFF_X al_4e658dcf (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[20]),
    .en(al_82faa065),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[20]));
  AL_DFF_X al_8e09f9d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[21]),
    .en(al_82faa065),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[21]));
  AL_DFF_X al_f0636598 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[22]),
    .en(al_82faa065),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[22]));
  AL_DFF_X al_806088f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[23]),
    .en(al_82faa065),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[23]));
  AL_DFF_X al_b244a282 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[24]),
    .en(al_82faa065),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[24]));
  AL_DFF_X al_e7214706 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[25]),
    .en(al_82faa065),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[25]));
  AL_DFF_X al_ca9bce13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[26]),
    .en(al_82faa065),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[26]));
  AL_DFF_X al_2009d0b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[27]),
    .en(al_82faa065),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[27]));
  AL_DFF_X al_e81fe6ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[28]),
    .en(al_82faa065),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[28]));
  AL_DFF_X al_94077685 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[2]),
    .en(al_82faa065),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[2]));
  AL_DFF_X al_5a9db3d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[29]),
    .en(al_82faa065),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[29]));
  AL_DFF_X al_f57b60e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[30]),
    .en(al_82faa065),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[30]));
  AL_DFF_X al_24f557ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[31]),
    .en(al_82faa065),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[31]));
  AL_DFF_X al_33016709 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[0]),
    .en(al_4965e5fa),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[32]));
  AL_DFF_X al_d9fd720b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[1]),
    .en(al_4965e5fa),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[33]));
  AL_DFF_X al_cff59033 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[2]),
    .en(al_4965e5fa),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[34]));
  AL_DFF_X al_36fd3bd3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[3]),
    .en(al_4965e5fa),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[35]));
  AL_DFF_X al_f1b05caf (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[4]),
    .en(al_4965e5fa),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[36]));
  AL_DFF_X al_df65b5da (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[5]),
    .en(al_4965e5fa),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[37]));
  AL_DFF_X al_25e82dde (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[6]),
    .en(al_4965e5fa),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[38]));
  AL_DFF_X al_e780f4d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[3]),
    .en(al_82faa065),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[3]));
  AL_DFF_X al_55e74ed7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[7]),
    .en(al_4965e5fa),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[39]));
  AL_DFF_X al_68770157 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[8]),
    .en(al_4965e5fa),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[40]));
  AL_DFF_X al_c338f8b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[9]),
    .en(al_4965e5fa),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[41]));
  AL_DFF_X al_de3ccacb (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[10]),
    .en(al_4965e5fa),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[42]));
  AL_DFF_X al_870b5695 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[11]),
    .en(al_4965e5fa),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[43]));
  AL_DFF_X al_d8c9a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[12]),
    .en(al_4965e5fa),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[44]));
  AL_DFF_X al_ffc85075 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[13]),
    .en(al_4965e5fa),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[45]));
  AL_DFF_X al_af9ce66a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[14]),
    .en(al_4965e5fa),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[46]));
  AL_DFF_X al_496bdce1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[15]),
    .en(al_4965e5fa),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[47]));
  AL_DFF_X al_f119555b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[16]),
    .en(al_4965e5fa),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[48]));
  AL_DFF_X al_ca953794 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[4]),
    .en(al_82faa065),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[4]));
  AL_DFF_X al_f711b2f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[17]),
    .en(al_4965e5fa),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[49]));
  AL_DFF_X al_853c2d30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[18]),
    .en(al_4965e5fa),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[50]));
  AL_DFF_X al_a7fe7c24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[19]),
    .en(al_4965e5fa),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[51]));
  AL_DFF_X al_8991048d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[20]),
    .en(al_4965e5fa),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[52]));
  AL_DFF_X al_a07a2ab5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[21]),
    .en(al_4965e5fa),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[53]));
  AL_DFF_X al_3decaa3c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[22]),
    .en(al_4965e5fa),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[54]));
  AL_DFF_X al_c0bbde78 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[23]),
    .en(al_4965e5fa),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[55]));
  AL_DFF_X al_eafd26b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[24]),
    .en(al_4965e5fa),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[56]));
  AL_DFF_X al_9ea33268 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[25]),
    .en(al_4965e5fa),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[57]));
  AL_DFF_X al_40980049 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[26]),
    .en(al_4965e5fa),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[58]));
  AL_DFF_X al_482e6132 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[5]),
    .en(al_82faa065),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[5]));
  AL_DFF_X al_21373840 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[27]),
    .en(al_4965e5fa),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[59]));
  AL_DFF_X al_9fece186 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[28]),
    .en(al_4965e5fa),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[60]));
  AL_DFF_X al_bf6675c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[29]),
    .en(al_4965e5fa),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[61]));
  AL_DFF_X al_e7d834ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[30]),
    .en(al_4965e5fa),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[62]));
  AL_DFF_X al_38f39387 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[31]),
    .en(al_4965e5fa),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[63]));
  AL_DFF_X al_6dffff0e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[6]),
    .en(al_82faa065),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[6]));
  AL_DFF_X al_235e2ea1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[7]),
    .en(al_82faa065),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[7]));
  AL_DFF_X al_cb24900c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[8]),
    .en(al_82faa065),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_d1b76c6b[8]));
  AL_DFF_X al_953bf09f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[0]));
  AL_DFF_X al_37f95a46 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[9]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[9]));
  AL_DFF_X al_72c867af (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[10]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[10]));
  AL_DFF_X al_585cfabe (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[11]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[11]));
  AL_DFF_X al_22691451 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[12]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[12]));
  AL_DFF_X al_e4fb78e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[13]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[13]));
  AL_DFF_X al_bad2054b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[14]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[14]));
  AL_DFF_X al_25aeff18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[15]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[15]));
  AL_DFF_X al_8852ca24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[16]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[16]));
  AL_DFF_X al_a4ad5075 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[17]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[17]));
  AL_DFF_X al_e3ecf00d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[18]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[18]));
  AL_DFF_X al_2f3593ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[1]));
  AL_DFF_X al_60c07466 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[19]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[19]));
  AL_DFF_X al_2176872c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[20]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[20]));
  AL_DFF_X al_6d82d94c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[21]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[21]));
  AL_DFF_X al_2fad62ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[22]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[22]));
  AL_DFF_X al_652499b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[23]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[23]));
  AL_DFF_X al_9df69309 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[24]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[24]));
  AL_DFF_X al_b07a3ff1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[25]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[25]));
  AL_DFF_X al_96269ff4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[26]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[26]));
  AL_DFF_X al_1bf6ab9e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[27]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[27]));
  AL_DFF_X al_2450e0a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[28]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[28]));
  AL_DFF_X al_aadf7880 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[2]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[2]));
  AL_DFF_X al_d2a185b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[29]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[29]));
  AL_DFF_X al_b633309b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[30]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[30]));
  AL_DFF_X al_cd181601 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[31]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[31]));
  AL_DFF_X al_f2772ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[32]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[32]));
  AL_DFF_X al_6ee2dc99 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[33]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[33]));
  AL_DFF_X al_82583a49 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[34]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[34]));
  AL_DFF_X al_d05026a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[35]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[35]));
  AL_DFF_X al_dbc6a958 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[36]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[36]));
  AL_DFF_X al_d22ea1e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[37]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[37]));
  AL_DFF_X al_d9f3e59a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[38]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[38]));
  AL_DFF_X al_79006f4f (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[3]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[3]));
  AL_DFF_X al_a643ae3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[39]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[39]));
  AL_DFF_X al_70ba7e23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[40]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[40]));
  AL_DFF_X al_742529f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[41]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[41]));
  AL_DFF_X al_2987796e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[42]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[42]));
  AL_DFF_X al_3577737c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[43]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[43]));
  AL_DFF_X al_3bb66476 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[44]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[44]));
  AL_DFF_X al_31d2684d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[45]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[45]));
  AL_DFF_X al_820a939d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[46]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[46]));
  AL_DFF_X al_c17314cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[47]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[47]));
  AL_DFF_X al_458bf6be (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[4]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[4]));
  AL_DFF_X al_16c19b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[5]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[5]));
  AL_DFF_X al_d6674ea9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[6]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[6]));
  AL_DFF_X al_426d1709 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[7]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[7]));
  AL_DFF_X al_c9748131 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_40f6174[8]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2408f449[8]));
  AL_DFF_X al_707ae6f3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[0]),
    .en(al_b7164eee),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[0]));
  AL_DFF_X al_11c5474f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[9]),
    .en(al_b7164eee),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[9]));
  AL_DFF_X al_68f57489 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[10]),
    .en(al_b7164eee),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[10]));
  AL_DFF_X al_c7cf5656 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[11]),
    .en(al_b7164eee),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[11]));
  AL_DFF_X al_a1e701e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[12]),
    .en(al_b7164eee),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[12]));
  AL_DFF_X al_47f08e9c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[13]),
    .en(al_b7164eee),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[13]));
  AL_DFF_X al_e594552b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[14]),
    .en(al_b7164eee),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[14]));
  AL_DFF_X al_d8f6be17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[15]),
    .en(al_b7164eee),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[15]));
  AL_DFF_X al_8c782e1b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[16]),
    .en(al_b7164eee),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[16]));
  AL_DFF_X al_2ea447f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[17]),
    .en(al_b7164eee),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[17]));
  AL_DFF_X al_994b49a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[18]),
    .en(al_b7164eee),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[18]));
  AL_DFF_X al_df828bec (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[1]),
    .en(al_b7164eee),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[1]));
  AL_DFF_X al_3a49df15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[19]),
    .en(al_b7164eee),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[19]));
  AL_DFF_X al_c20edec8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[20]),
    .en(al_b7164eee),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[20]));
  AL_DFF_X al_a5c1101b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[21]),
    .en(al_b7164eee),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[21]));
  AL_DFF_X al_b9cd7639 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[22]),
    .en(al_b7164eee),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[22]));
  AL_DFF_X al_ca06c2b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[23]),
    .en(al_b7164eee),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[23]));
  AL_DFF_X al_781b9488 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[24]),
    .en(al_b7164eee),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[24]));
  AL_DFF_X al_e4ee15fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[25]),
    .en(al_b7164eee),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[25]));
  AL_DFF_X al_165feba1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[26]),
    .en(al_b7164eee),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[26]));
  AL_DFF_X al_6cb9c9a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[27]),
    .en(al_b7164eee),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[27]));
  AL_DFF_X al_aa4939cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[28]),
    .en(al_b7164eee),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[28]));
  AL_DFF_X al_287b5ca6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[2]),
    .en(al_b7164eee),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[2]));
  AL_DFF_X al_f10e5916 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[29]),
    .en(al_b7164eee),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[29]));
  AL_DFF_X al_b02933e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[30]),
    .en(al_b7164eee),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[30]));
  AL_DFF_X al_90abb62d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[31]),
    .en(al_b7164eee),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[31]));
  AL_DFF_X al_30acd42b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[0]),
    .en(al_e3838f69),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[32]));
  AL_DFF_X al_5e02a189 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[1]),
    .en(al_e3838f69),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[33]));
  AL_DFF_X al_e1731a97 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[2]),
    .en(al_e3838f69),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[34]));
  AL_DFF_X al_deccbb34 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[3]),
    .en(al_e3838f69),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[35]));
  AL_DFF_X al_44140212 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[4]),
    .en(al_e3838f69),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[36]));
  AL_DFF_X al_4e8d120c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[5]),
    .en(al_e3838f69),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[37]));
  AL_DFF_X al_a3c9cf25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[6]),
    .en(al_e3838f69),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[38]));
  AL_DFF_X al_a5e82312 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[3]),
    .en(al_b7164eee),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[3]));
  AL_DFF_X al_db73abf8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[7]),
    .en(al_e3838f69),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[39]));
  AL_DFF_X al_d39898cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[8]),
    .en(al_e3838f69),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[40]));
  AL_DFF_X al_86fe0328 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[9]),
    .en(al_e3838f69),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[41]));
  AL_DFF_X al_64af99fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[10]),
    .en(al_e3838f69),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[42]));
  AL_DFF_X al_7fba60db (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[11]),
    .en(al_e3838f69),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[43]));
  AL_DFF_X al_5b4866b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[12]),
    .en(al_e3838f69),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[44]));
  AL_DFF_X al_649a52f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[13]),
    .en(al_e3838f69),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[45]));
  AL_DFF_X al_123bea8e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[14]),
    .en(al_e3838f69),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[46]));
  AL_DFF_X al_d446d779 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[15]),
    .en(al_e3838f69),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[47]));
  AL_DFF_X al_c8580d45 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[16]),
    .en(al_e3838f69),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[48]));
  AL_DFF_X al_61552569 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[4]),
    .en(al_b7164eee),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[4]));
  AL_DFF_X al_69da2544 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[17]),
    .en(al_e3838f69),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[49]));
  AL_DFF_X al_33f7bdab (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[18]),
    .en(al_e3838f69),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[50]));
  AL_DFF_X al_bf59d3c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[19]),
    .en(al_e3838f69),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[51]));
  AL_DFF_X al_dad3eaf0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[20]),
    .en(al_e3838f69),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[52]));
  AL_DFF_X al_7e800419 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[21]),
    .en(al_e3838f69),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[53]));
  AL_DFF_X al_6d962d81 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[22]),
    .en(al_e3838f69),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[54]));
  AL_DFF_X al_9e2505d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[23]),
    .en(al_e3838f69),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[55]));
  AL_DFF_X al_b2564d86 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[24]),
    .en(al_e3838f69),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[56]));
  AL_DFF_X al_10993021 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[25]),
    .en(al_e3838f69),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[57]));
  AL_DFF_X al_e7085f15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[26]),
    .en(al_e3838f69),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[58]));
  AL_DFF_X al_8a34dba7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[5]),
    .en(al_b7164eee),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[5]));
  AL_DFF_X al_9a18df65 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[27]),
    .en(al_e3838f69),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[59]));
  AL_DFF_X al_a3d8173a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[28]),
    .en(al_e3838f69),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[60]));
  AL_DFF_X al_7bda8ba8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[29]),
    .en(al_e3838f69),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[61]));
  AL_DFF_X al_3f9147bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[30]),
    .en(al_e3838f69),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[62]));
  AL_DFF_X al_85932db0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[31]),
    .en(al_e3838f69),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[63]));
  AL_DFF_X al_c5ff4e47 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[6]),
    .en(al_b7164eee),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[6]));
  AL_DFF_X al_40c54362 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[7]),
    .en(al_b7164eee),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[7]));
  AL_DFF_X al_d886c61d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(s_axi_wdata[8]),
    .en(al_b7164eee),
    .sr(al_81344cef),
    .ss(1'b0),
    .q(al_752f7592[8]));
  AL_DFF_X al_659c5183 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_6aaeddf4),
    .d(al_e6b493f[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a4fb2b45));
  AL_DFF_X al_335a39b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_6aaeddf4),
    .d(al_e6b493f[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a6bba48));
  AL_DFF_X al_34c270b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_6aaeddf4),
    .d(al_e6b493f[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c3e9514));
  AL_DFF_X al_80f5cace (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_6aaeddf4),
    .d(al_e6b493f[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1396ae3));
  AL_DFF_X al_c026dbd1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_6aaeddf4),
    .d(al_e6b493f[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_da9f8ded));
  AL_DFF_X al_8a219ef8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_6aaeddf4),
    .d(al_e6b493f[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_655153ec));
  AL_DFF_X al_aeb24fc9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_6aaeddf4),
    .d(al_e6b493f[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ba02654));
  AL_DFF_X al_24b9abf6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_6aaeddf4),
    .d(al_e6b493f[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9993ad5e));
  AL_DFF_X al_cff971f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_6aaeddf4),
    .d(al_e6b493f[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29e11b90));
  AL_DFF_X al_64280ddf (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_6aaeddf4),
    .d(al_e6b493f[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a1cb58));
  AL_DFF_X al_e409aef3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_6aaeddf4),
    .d(al_e6b493f[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_989215e7));
  AL_DFF_X al_d0cc875 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_6aaeddf4),
    .d(al_e6b493f[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac9336a));
  AL_DFF_X al_8891cbd9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_6aaeddf4),
    .d(al_e6b493f[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c616a92));
  AL_DFF_X al_970233a (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_6aaeddf4),
    .d(al_e6b493f[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e19dcc16));
  AL_DFF_X al_4da61663 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_6aaeddf4),
    .d(al_e6b493f[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a4c57dd8));
  AL_DFF_X al_96449dd7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_6aaeddf4),
    .d(al_e6b493f[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4b485d4));
  AL_DFF_X al_7fe63eb9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_6aaeddf4),
    .d(al_e6b493f[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a880ef2c));
  AL_DFF_X al_fabba4d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_6aaeddf4),
    .d(al_e6b493f[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1974d963));
  AL_DFF_X al_243584ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_6aaeddf4),
    .d(al_e6b493f[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b3009928));
  AL_DFF_X al_21ba7078 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_6aaeddf4),
    .d(al_e6b493f[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f13bd74f));
  AL_DFF_X al_c43dd0fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_6aaeddf4),
    .d(al_e6b493f[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ad06c7e));
  AL_DFF_X al_e072813a (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_6aaeddf4),
    .d(al_e6b493f[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_159c9d41));
  AL_DFF_X al_3b8fd63e (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_6aaeddf4),
    .d(al_e6b493f[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fefd5fd3));
  AL_DFF_X al_6f18e988 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_6aaeddf4),
    .d(al_e6b493f[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ca969cfa));
  AL_DFF_X al_70423b07 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_6aaeddf4),
    .d(al_e6b493f[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_dd993167));
  AL_DFF_X al_d636ea75 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_6aaeddf4),
    .d(al_e6b493f[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4285f2d3));
  AL_DFF_X al_6594dd98 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_6aaeddf4),
    .d(al_e6b493f[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8b78b709));
  AL_DFF_X al_79e72508 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_6aaeddf4),
    .d(al_e6b493f[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c40403fa));
  AL_DFF_X al_213f7ae6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_6aaeddf4),
    .d(al_e6b493f[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6be24f));
  AL_DFF_X al_103999f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_6aaeddf4),
    .d(al_e6b493f[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad7719c4));
  AL_DFF_X al_4d90bc51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_6aaeddf4),
    .d(al_e6b493f[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_eaf2c767));
  AL_DFF_X al_815167ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(~al_6aaeddf4),
    .d(al_e6b493f[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8b492536));
  AL_DFF_X al_60e40fe6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[0]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[0]));
  AL_DFF_X al_44dba831 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[9]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[9]));
  AL_DFF_X al_e4c08a39 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[10]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[10]));
  AL_DFF_X al_7e629447 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[11]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[11]));
  AL_DFF_X al_5427dc42 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[12]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[12]));
  AL_DFF_X al_33cc04e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[13]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[13]));
  AL_DFF_X al_798ec84b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[14]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[14]));
  AL_DFF_X al_e3299273 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[15]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[15]));
  AL_DFF_X al_4bc6b914 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[16]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[16]));
  AL_DFF_X al_2c101db6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[17]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[17]));
  AL_DFF_X al_202962f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[18]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[18]));
  AL_DFF_X al_f15b8e07 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[1]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[1]));
  AL_DFF_X al_12f13fa5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[19]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[19]));
  AL_DFF_X al_5ec0d63 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[20]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[20]));
  AL_DFF_X al_c2067d51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[21]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[21]));
  AL_DFF_X al_5f19ff7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[22]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[22]));
  AL_DFF_X al_67891e13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[23]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[23]));
  AL_DFF_X al_3cf90f0d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[24]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[24]));
  AL_DFF_X al_175ca01 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[25]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[25]));
  AL_DFF_X al_485cc5fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[26]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[26]));
  AL_DFF_X al_5b277c0a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[27]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[27]));
  AL_DFF_X al_403972d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[28]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[28]));
  AL_DFF_X al_16ef1bc6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[2]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[2]));
  AL_DFF_X al_4c92ea47 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[29]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[29]));
  AL_DFF_X al_1d254ffd (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[30]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[30]));
  AL_DFF_X al_5d2f7bc7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[31]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[31]));
  AL_DFF_X al_9a903262 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[32]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[32]));
  AL_DFF_X al_66e6d68d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[33]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[33]));
  AL_DFF_X al_2cbd5ddc (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[34]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[34]));
  AL_DFF_X al_c91766c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[35]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[35]));
  AL_DFF_X al_7c99a03b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[36]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[36]));
  AL_DFF_X al_f3c55d31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[37]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[37]));
  AL_DFF_X al_e02bb120 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[38]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[38]));
  AL_DFF_X al_46094d5e (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[3]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[3]));
  AL_DFF_X al_5df11b4a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[39]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[39]));
  AL_DFF_X al_e2b2ebf2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[40]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[40]));
  AL_DFF_X al_8c2f5f2d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[41]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[41]));
  AL_DFF_X al_b191982a (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[42]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[42]));
  AL_DFF_X al_1bdc6fe1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[43]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[43]));
  AL_DFF_X al_5b259a9c (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[44]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[44]));
  AL_DFF_X al_d10721e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[45]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[45]));
  AL_DFF_X al_9e2a5d83 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[46]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[46]));
  AL_DFF_X al_656af615 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[47]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[47]));
  AL_DFF_X al_40acceaa (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[4]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[4]));
  AL_DFF_X al_15305606 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[5]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[5]));
  AL_DFF_X al_fa6c9597 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[6]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[6]));
  AL_DFF_X al_91fa8105 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[7]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[7]));
  AL_DFF_X al_50abd803 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_f0cac652[8]),
    .en(rx_clk_en),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2bdcc449[8]));
  AL_DFF_X al_a16cf221 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[0]));
  AL_DFF_X al_25cc6963 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[9]));
  AL_DFF_X al_e976fac2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[10]));
  AL_DFF_X al_bbf2608e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[11]));
  AL_DFF_X al_4573fbba (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[12]));
  AL_DFF_X al_367e2412 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[13]));
  AL_DFF_X al_6519478 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[14]));
  AL_DFF_X al_e86d906b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[15]));
  AL_DFF_X al_d3d20149 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[16]));
  AL_DFF_X al_996e854c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[17]));
  AL_DFF_X al_bd227e8b (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[18]));
  AL_DFF_X al_4b642686 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[1]));
  AL_DFF_X al_73b6e493 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[19]));
  AL_DFF_X al_5de2c6ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[20]));
  AL_DFF_X al_76af1bad (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[21]));
  AL_DFF_X al_3d6f9cfc (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[22]));
  AL_DFF_X al_a4490d70 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[23]));
  AL_DFF_X al_caa47320 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[24]));
  AL_DFF_X al_dc73db1a (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[25]));
  AL_DFF_X al_c2bbc83c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[26]));
  AL_DFF_X al_12e272e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[27]));
  AL_DFF_X al_4390f4e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[28]));
  AL_DFF_X al_8a19c0c (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[2]));
  AL_DFF_X al_2c055775 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[29]));
  AL_DFF_X al_25b08a88 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[30]));
  AL_DFF_X al_e9f6ab25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[31]));
  AL_DFF_X al_8e8f78bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[32]));
  AL_DFF_X al_a9ab2895 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[33]));
  AL_DFF_X al_96b7734e (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[34]));
  AL_DFF_X al_8ed062b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[35]));
  AL_DFF_X al_c4bdeede (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[36]));
  AL_DFF_X al_fd3fdbc8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[37]));
  AL_DFF_X al_c19aa374 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[38]));
  AL_DFF_X al_f19ef88f (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[3]));
  AL_DFF_X al_663bd4c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[39]));
  AL_DFF_X al_af0193a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[40]));
  AL_DFF_X al_7ff01e2d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[41]));
  AL_DFF_X al_2c4007f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[42]));
  AL_DFF_X al_3f1bbe0d (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[43]));
  AL_DFF_X al_68c15bf5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[44]));
  AL_DFF_X al_a51abd68 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[45]));
  AL_DFF_X al_76bee1c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[46]));
  AL_DFF_X al_4d61d568 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[47]));
  AL_DFF_X al_a826fb12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[4]));
  AL_DFF_X al_51f9d165 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[5]));
  AL_DFF_X al_7c582a46 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[6]));
  AL_DFF_X al_5469e65 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[7]));
  AL_DFF_X al_bdca02d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_9db0b0fa[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_49a90ce2[8]));
  AL_DFF_X al_22be2317 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_f3e1aff9),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b9297703[0]));
  AL_DFF_X al_2a1693a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_10307540),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b9297703[1]));
  AL_MAP_LUT6 #(
    .EQN("(F*E*~D*~C*~B*A)"),
    .INIT(64'h0002000000000000))
    al_6cdb7d4e (
    .a(s_axi_awaddr[7]),
    .b(s_axi_awaddr[6]),
    .c(s_axi_awaddr[5]),
    .d(s_axi_awaddr[4]),
    .e(s_axi_awvalid),
    .f(s_axi_wvalid),
    .o(al_a53ff9fc));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*C*~B*A)"),
    .INIT(32'h00002000))
    al_6344a784 (
    .a(al_a53ff9fc),
    .b(s_axi_awaddr[3]),
    .c(s_axi_awaddr[2]),
    .d(s_axi_awaddr[1]),
    .e(s_axi_awaddr[0]),
    .o(al_dc8505e1));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'h0d08))
    al_82d746d8 (
    .a(al_dc8505e1),
    .b(s_axi_wdata[16]),
    .c(al_81344cef),
    .d(al_b9297703[0]),
    .o(al_f3e1aff9));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'h0d08))
    al_6069dd8b (
    .a(al_dc8505e1),
    .b(s_axi_wdata[19]),
    .c(al_81344cef),
    .d(al_b9297703[3]),
    .o(al_bfa502a9));
  AL_DFF_X al_94d4e092 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_332cacdd),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b9297703[2]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'h0d08))
    al_282efd84 (
    .a(al_dc8505e1),
    .b(s_axi_wdata[18]),
    .c(al_81344cef),
    .d(al_b9297703[2]),
    .o(al_332cacdd));
  AL_MAP_LUT4 #(
    .EQN("(~C*(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'h0d08))
    al_c0e4943e (
    .a(al_dc8505e1),
    .b(s_axi_wdata[17]),
    .c(al_81344cef),
    .d(al_b9297703[1]),
    .o(al_10307540));
  AL_DFF_X al_534d8541 (
    .ar(1'b0),
    .as(1'b0),
    .clk(s_axi_aclk),
    .d(al_bfa502a9),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b9297703[3]));
  AL_DFF_X al_4344e99d (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_ecfcb422[3]),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(rx_status_vector[4]));
  AL_DFF_X al_84dcc17b (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_6ab23518),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_3edda74b));
  AL_MAP_LUT3 #(
    .EQN("(~A*~B*~C+A*~B*C)"),
    .INIT(8'b00100001))
    al_8125417f (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_d0555e9d[2]),
    .o(al_5fe249d5[0]));
  AL_MAP_LUT3 #(
    .EQN("(A*~B*~C+~A*B*~C)"),
    .INIT(8'b00000110))
    al_a792efda (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .c(al_d0555e9d[2]),
    .o(al_5fe249d5[7]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_93bb2ed7 (
    .a(al_d0555e9d[0]),
    .b(al_d0555e9d[1]),
    .o(al_968fd17c));
  AL_MAP_LUT6 #(
    .EQN("(~D*~C*~B*~A*~(F@E))"),
    .INIT(64'h0001000000000001))
    al_eb52d69d (
    .a(al_e8c5f626[2]),
    .b(al_e8c5f626[3]),
    .c(al_e8c5f626[4]),
    .d(al_e8c5f626[5]),
    .e(al_e8c5f626[7]),
    .f(al_5fe249d5[7]),
    .o(al_4f2f7ae3));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*A))"),
    .INIT(8'h0d))
    al_416ca6ba (
    .a(al_132ae268),
    .b(al_30b5e311),
    .c(al_3edda74b),
    .o(al_904a5dce));
  AL_MAP_LUT5 #(
    .EQN("(~A*(~(C)*~(D)*~((~E*B))+C*D*(~E*B)))"),
    .INIT(32'h00054001))
    al_f1d5615 (
    .a(al_904a5dce),
    .b(al_968fd17c),
    .c(al_e8c5f626[1]),
    .d(al_e8c5f626[6]),
    .e(al_d0555e9d[2]),
    .o(al_fc8b055a));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    al_e4fe7361 (
    .a(al_fc8b055a),
    .b(al_4f2f7ae3),
    .c(al_e8c5f626[0]),
    .d(al_5fe249d5[0]),
    .o(al_6ab23518));
  AL_DFF_X al_3bcccf83 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_1bc55ab2),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_8399b753));
  AL_DFF_X al_f1e68919 (
    .ar(1'b0),
    .as(1'b0),
    .clk(rx_mac_clk),
    .d(al_3e178366),
    .en(rx_clk_en),
    .sr(al_ff9a7266),
    .ss(1'b0),
    .q(al_536b4576));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_fa020be7 (
    .a(al_25215c55[0]),
    .b(al_25215c55[1]),
    .o(al_72f5321b));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_53c015fe (
    .a(al_6b181c0),
    .b(al_7968b2a5),
    .o(mdio_clk));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_979c3f3f (
    .a(al_abc98a52),
    .b(al_678e4333),
    .c(al_8b780845),
    .o(al_6de80447));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_c35e3378 (
    .a(al_6de80447),
    .b(al_1feb4c09),
    .o(rx_status_vector[23]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_3be2914f (
    .a(al_2bb2d81d),
    .b(al_1feb4c09),
    .c(al_8e811a01),
    .o(rx_status_vector[24]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_e9858ef3 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[0]),
    .d(al_d1b76c6b[0]),
    .e(al_752f7592[0]),
    .o(al_810ba8de));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_8c397c3f (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[32]),
    .d(al_d1b76c6b[32]),
    .e(al_752f7592[32]),
    .o(al_8b51ab4));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_9f16686c (
    .a(al_175588ec),
    .b(al_8b51ab4),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_b9297703[2]),
    .f(al_b9297703[3]),
    .o(al_f8a9808f));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))"),
    .INIT(32'h22200200))
    al_d8aec332 (
    .a(al_175588ec),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_49a90ce2[0]),
    .e(al_49a90ce2[32]),
    .o(al_2da9429f));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_162714cb (
    .a(al_fc03cb77),
    .b(al_f8a9808f),
    .c(al_2da9429f),
    .d(al_810ba8de),
    .e(al_88fb5330[0]),
    .f(al_a9336f5),
    .o(al_e6b493f[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_d960c7a7 (
    .a(al_e6b493f[0]),
    .b(al_6aaeddf4),
    .c(al_e4b485d4),
    .o(s_axi_rdata[0]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_9d8f26d9 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[10]),
    .d(al_d1b76c6b[10]),
    .e(al_752f7592[10]),
    .o(al_1d01387));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_9513daa3 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[42]),
    .d(al_d1b76c6b[42]),
    .e(al_752f7592[42]),
    .o(al_8e145c1c));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_80339ef1 (
    .a(al_175588ec),
    .b(al_8e145c1c),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_b9297703[2]),
    .f(al_b9297703[3]),
    .o(al_c9f27122));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))"),
    .INIT(32'h22200200))
    al_d3917c52 (
    .a(al_175588ec),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_49a90ce2[10]),
    .e(al_49a90ce2[42]),
    .o(al_f5bbf69e));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_89b3ed75 (
    .a(al_fc03cb77),
    .b(al_c9f27122),
    .c(al_f5bbf69e),
    .d(al_1d01387),
    .e(al_88fb5330[10]),
    .f(al_a9336f5),
    .o(al_e6b493f[10]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_932ea8d8 (
    .a(al_e6b493f[10]),
    .b(al_6aaeddf4),
    .c(al_4285f2d3),
    .o(s_axi_rdata[10]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_8935f2cd (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[11]),
    .d(al_d1b76c6b[11]),
    .e(al_752f7592[11]),
    .o(al_1caff122));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_d7fbaccd (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[43]),
    .d(al_d1b76c6b[43]),
    .e(al_752f7592[43]),
    .o(al_826fce19));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_ed1d54d8 (
    .a(al_175588ec),
    .b(al_826fce19),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_b9297703[2]),
    .f(al_b9297703[3]),
    .o(al_3a099803));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))"),
    .INIT(32'h22200200))
    al_beba8616 (
    .a(al_175588ec),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_49a90ce2[11]),
    .e(al_49a90ce2[43]),
    .o(al_a8b162ca));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_62af4930 (
    .a(al_fc03cb77),
    .b(al_3a099803),
    .c(al_a8b162ca),
    .d(al_1caff122),
    .e(al_88fb5330[11]),
    .f(al_a9336f5),
    .o(al_e6b493f[11]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_8e952a89 (
    .a(al_e6b493f[11]),
    .b(al_6aaeddf4),
    .c(al_8b78b709),
    .o(s_axi_rdata[11]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_760683d5 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[12]),
    .d(al_d1b76c6b[12]),
    .e(al_752f7592[12]),
    .o(al_acabe8fb));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_652169a1 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[44]),
    .d(al_d1b76c6b[44]),
    .e(al_752f7592[44]),
    .o(al_46ece34d));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_48b1bf9e (
    .a(al_175588ec),
    .b(al_46ece34d),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_b9297703[2]),
    .f(al_b9297703[3]),
    .o(al_1d49aa78));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))"),
    .INIT(32'h22200200))
    al_86c9f18f (
    .a(al_175588ec),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_49a90ce2[12]),
    .e(al_49a90ce2[44]),
    .o(al_f474e268));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_9e4693c2 (
    .a(al_fc03cb77),
    .b(al_1d49aa78),
    .c(al_f474e268),
    .d(al_acabe8fb),
    .e(al_88fb5330[12]),
    .f(al_a9336f5),
    .o(al_e6b493f[12]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_952ddb35 (
    .a(al_e6b493f[12]),
    .b(al_6aaeddf4),
    .c(al_c40403fa),
    .o(s_axi_rdata[12]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_95243338 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[13]),
    .d(al_d1b76c6b[13]),
    .e(al_752f7592[13]),
    .o(al_9fcf7528));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_c955b043 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[45]),
    .d(al_d1b76c6b[45]),
    .e(al_752f7592[45]),
    .o(al_4beb6793));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_f310fe51 (
    .a(al_175588ec),
    .b(al_4beb6793),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_b9297703[2]),
    .f(al_b9297703[3]),
    .o(al_67882c63));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))"),
    .INIT(32'h22200200))
    al_b290fe81 (
    .a(al_175588ec),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_49a90ce2[13]),
    .e(al_49a90ce2[45]),
    .o(al_8952b398));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_32ba3cda (
    .a(al_fc03cb77),
    .b(al_67882c63),
    .c(al_8952b398),
    .d(al_9fcf7528),
    .e(al_88fb5330[13]),
    .f(al_a9336f5),
    .o(al_e6b493f[13]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_e8487bc4 (
    .a(al_e6b493f[13]),
    .b(al_6aaeddf4),
    .c(al_b6be24f),
    .o(s_axi_rdata[13]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_8c5df2fe (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[14]),
    .d(al_d1b76c6b[14]),
    .e(al_752f7592[14]),
    .o(al_5006fa3b));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_f5cf77c1 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[46]),
    .d(al_d1b76c6b[46]),
    .e(al_752f7592[46]),
    .o(al_53f52d8d));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_62df8762 (
    .a(al_175588ec),
    .b(al_53f52d8d),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_b9297703[2]),
    .f(al_b9297703[3]),
    .o(al_133f55a2));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))"),
    .INIT(32'h22200200))
    al_79374e07 (
    .a(al_175588ec),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_49a90ce2[14]),
    .e(al_49a90ce2[46]),
    .o(al_78512832));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_c7f66efb (
    .a(al_fc03cb77),
    .b(al_133f55a2),
    .c(al_78512832),
    .d(al_5006fa3b),
    .e(al_88fb5330[14]),
    .f(al_a9336f5),
    .o(al_e6b493f[14]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_b1aa3a41 (
    .a(al_e6b493f[14]),
    .b(al_6aaeddf4),
    .c(al_ad7719c4),
    .o(s_axi_rdata[14]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_356e2313 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[15]),
    .d(al_d1b76c6b[15]),
    .e(al_752f7592[15]),
    .o(al_9fbaf8f2));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_70e4251c (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[47]),
    .d(al_d1b76c6b[47]),
    .e(al_752f7592[47]),
    .o(al_dbb71724));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_22cf0863 (
    .a(al_175588ec),
    .b(al_dbb71724),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_b9297703[2]),
    .f(al_b9297703[3]),
    .o(al_d849110a));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))"),
    .INIT(32'h22200200))
    al_85892546 (
    .a(al_175588ec),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_49a90ce2[15]),
    .e(al_49a90ce2[47]),
    .o(al_715827e7));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_e87298d (
    .a(al_fc03cb77),
    .b(al_d849110a),
    .c(al_715827e7),
    .d(al_9fbaf8f2),
    .e(al_88fb5330[15]),
    .f(al_a9336f5),
    .o(al_e6b493f[15]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_728122bd (
    .a(al_e6b493f[15]),
    .b(al_6aaeddf4),
    .c(al_eaf2c767),
    .o(s_axi_rdata[15]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_2d31bc8d (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[16]),
    .d(al_d1b76c6b[16]),
    .e(al_752f7592[16]),
    .o(al_18c1e35a));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_19d6b37c (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[48]),
    .d(al_d1b76c6b[48]),
    .e(al_752f7592[48]),
    .o(al_662270e8));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(~D*B)*~(~E*A))"),
    .INIT(64'h0f030501ff335511))
    al_8dcd45c9 (
    .a(al_627de329),
    .b(al_fc03cb77),
    .c(al_ce826c89),
    .d(al_18c1e35a),
    .e(al_662270e8),
    .f(al_49a90ce2[16]),
    .o(al_a03de72f));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))*~(B)+~E*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*~(B)+~(~E)*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*B+~E*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*B)"),
    .INIT(32'h77f344c0))
    al_1c830f5d (
    .a(al_a03de72f),
    .b(al_6aaeddf4),
    .c(al_88fb5330[16]),
    .d(al_a9336f5),
    .e(al_8b492536),
    .o(s_axi_rdata[16]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_a7082b37 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[17]),
    .d(al_d1b76c6b[17]),
    .e(al_752f7592[17]),
    .o(al_42966d4a));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_93d562e5 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[49]),
    .d(al_d1b76c6b[49]),
    .e(al_752f7592[49]),
    .o(al_8c6ac38c));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(~D*B)*~(~E*A))"),
    .INIT(64'h0f030501ff335511))
    al_65fe8947 (
    .a(al_627de329),
    .b(al_fc03cb77),
    .c(al_ce826c89),
    .d(al_42966d4a),
    .e(al_8c6ac38c),
    .f(al_49a90ce2[17]),
    .o(al_81681eb));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))*~(B)+~E*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*~(B)+~(~E)*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*B+~E*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*B)"),
    .INIT(32'h77f344c0))
    al_a3679761 (
    .a(al_81681eb),
    .b(al_6aaeddf4),
    .c(al_88fb5330[17]),
    .d(al_a9336f5),
    .e(al_a4fb2b45),
    .o(s_axi_rdata[17]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_ff9ff38e (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[18]),
    .d(al_d1b76c6b[18]),
    .e(al_752f7592[18]),
    .o(al_3aae9c28));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_21461c20 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[50]),
    .d(al_d1b76c6b[50]),
    .e(al_752f7592[50]),
    .o(al_346eaec2));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(~D*B)*~(~E*A))"),
    .INIT(64'h0f030501ff335511))
    al_393de1b4 (
    .a(al_627de329),
    .b(al_fc03cb77),
    .c(al_ce826c89),
    .d(al_3aae9c28),
    .e(al_346eaec2),
    .f(al_49a90ce2[18]),
    .o(al_644f021d));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))*~(B)+~E*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*~(B)+~(~E)*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*B+~E*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*B)"),
    .INIT(32'h77f344c0))
    al_f1e7f594 (
    .a(al_644f021d),
    .b(al_6aaeddf4),
    .c(al_88fb5330[18]),
    .d(al_a9336f5),
    .e(al_6a6bba48),
    .o(s_axi_rdata[18]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_fe8ea8ec (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[19]),
    .d(al_d1b76c6b[19]),
    .e(al_752f7592[19]),
    .o(al_be16aa76));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_333eb66e (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[51]),
    .d(al_d1b76c6b[51]),
    .e(al_752f7592[51]),
    .o(al_b2b8b63f));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(~D*B)*~(~E*A))"),
    .INIT(64'h0f030501ff335511))
    al_8143caa4 (
    .a(al_627de329),
    .b(al_fc03cb77),
    .c(al_ce826c89),
    .d(al_be16aa76),
    .e(al_b2b8b63f),
    .f(al_49a90ce2[19]),
    .o(al_f4252f15));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))*~(B)+~E*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*~(B)+~(~E)*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*B+~E*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*B)"),
    .INIT(32'h77f344c0))
    al_4ffe8138 (
    .a(al_f4252f15),
    .b(al_6aaeddf4),
    .c(al_88fb5330[19]),
    .d(al_a9336f5),
    .e(al_c3e9514),
    .o(s_axi_rdata[19]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_a95349da (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[1]),
    .d(al_d1b76c6b[1]),
    .e(al_752f7592[1]),
    .o(al_5fd6768b));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_964b914f (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[33]),
    .d(al_d1b76c6b[33]),
    .e(al_752f7592[33]),
    .o(al_38ea72f1));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_4705734b (
    .a(al_175588ec),
    .b(al_38ea72f1),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_b9297703[2]),
    .f(al_b9297703[3]),
    .o(al_50c6f567));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))"),
    .INIT(32'h22200200))
    al_911365c7 (
    .a(al_175588ec),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_49a90ce2[1]),
    .e(al_49a90ce2[33]),
    .o(al_64bc3920));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_690c493d (
    .a(al_fc03cb77),
    .b(al_50c6f567),
    .c(al_64bc3920),
    .d(al_5fd6768b),
    .e(al_88fb5330[1]),
    .f(al_a9336f5),
    .o(al_e6b493f[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_e76f55f7 (
    .a(al_e6b493f[1]),
    .b(al_6aaeddf4),
    .c(al_a880ef2c),
    .o(s_axi_rdata[1]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_ef452774 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[20]),
    .d(al_d1b76c6b[20]),
    .e(al_752f7592[20]),
    .o(al_ac5af120));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_906fd266 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[52]),
    .d(al_d1b76c6b[52]),
    .e(al_752f7592[52]),
    .o(al_d9170e3));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(~D*B)*~(~E*A))"),
    .INIT(64'h0f030501ff335511))
    al_fa16511d (
    .a(al_627de329),
    .b(al_fc03cb77),
    .c(al_ce826c89),
    .d(al_ac5af120),
    .e(al_d9170e3),
    .f(al_49a90ce2[20]),
    .o(al_61fb0a6));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))*~(B)+~E*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*~(B)+~(~E)*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*B+~E*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*B)"),
    .INIT(32'h77f344c0))
    al_cd791c67 (
    .a(al_61fb0a6),
    .b(al_6aaeddf4),
    .c(al_88fb5330[20]),
    .d(al_a9336f5),
    .e(al_f1396ae3),
    .o(s_axi_rdata[20]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_5ea1e60b (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[21]),
    .d(al_d1b76c6b[21]),
    .e(al_752f7592[21]),
    .o(al_41b2f611));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_dca24c8f (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[53]),
    .d(al_d1b76c6b[53]),
    .e(al_752f7592[53]),
    .o(al_d7707346));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(~D*B)*~(~E*A))"),
    .INIT(64'h0f030501ff335511))
    al_afb7c2d5 (
    .a(al_627de329),
    .b(al_fc03cb77),
    .c(al_ce826c89),
    .d(al_41b2f611),
    .e(al_d7707346),
    .f(al_49a90ce2[21]),
    .o(al_3b505c23));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))*~(B)+~E*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*~(B)+~(~E)*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*B+~E*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*B)"),
    .INIT(32'h77f344c0))
    al_f7550574 (
    .a(al_3b505c23),
    .b(al_6aaeddf4),
    .c(al_88fb5330[21]),
    .d(al_a9336f5),
    .e(al_da9f8ded),
    .o(s_axi_rdata[21]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_496e42c5 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[22]),
    .d(al_d1b76c6b[22]),
    .e(al_752f7592[22]),
    .o(al_127a14bf));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_dc8f9434 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[54]),
    .d(al_d1b76c6b[54]),
    .e(al_752f7592[54]),
    .o(al_4dd161f2));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(~D*B)*~(~E*A))"),
    .INIT(64'h0f030501ff335511))
    al_c866ca5 (
    .a(al_627de329),
    .b(al_fc03cb77),
    .c(al_ce826c89),
    .d(al_127a14bf),
    .e(al_4dd161f2),
    .f(al_49a90ce2[22]),
    .o(al_179835d0));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))*~(B)+~E*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*~(B)+~(~E)*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*B+~E*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*B)"),
    .INIT(32'h77f344c0))
    al_4965d6d6 (
    .a(al_179835d0),
    .b(al_6aaeddf4),
    .c(al_88fb5330[22]),
    .d(al_a9336f5),
    .e(al_655153ec),
    .o(s_axi_rdata[22]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_12727fd8 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[23]),
    .d(al_d1b76c6b[23]),
    .e(al_752f7592[23]),
    .o(al_8f322b4));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_2a17bbdb (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[55]),
    .d(al_d1b76c6b[55]),
    .e(al_752f7592[55]),
    .o(al_11c159a));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(~D*B)*~(~E*A))"),
    .INIT(64'h0f030501ff335511))
    al_fb24d746 (
    .a(al_627de329),
    .b(al_fc03cb77),
    .c(al_ce826c89),
    .d(al_8f322b4),
    .e(al_11c159a),
    .f(al_49a90ce2[23]),
    .o(al_7cd2fee3));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))*~(B)+~E*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*~(B)+~(~E)*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*B+~E*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*B)"),
    .INIT(32'h77f344c0))
    al_d3763c57 (
    .a(al_7cd2fee3),
    .b(al_6aaeddf4),
    .c(al_88fb5330[23]),
    .d(al_a9336f5),
    .e(al_8ba02654),
    .o(s_axi_rdata[23]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_12bae85f (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[24]),
    .d(al_d1b76c6b[24]),
    .e(al_752f7592[24]),
    .o(al_64d29977));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_2526ac3b (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[56]),
    .d(al_d1b76c6b[56]),
    .e(al_752f7592[56]),
    .o(al_609ad6f2));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(~D*B)*~(~E*A))"),
    .INIT(64'h0f030501ff335511))
    al_2f5523e9 (
    .a(al_627de329),
    .b(al_fc03cb77),
    .c(al_ce826c89),
    .d(al_64d29977),
    .e(al_609ad6f2),
    .f(al_49a90ce2[24]),
    .o(al_70727c2f));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))*~(B)+~E*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*~(B)+~(~E)*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*B+~E*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*B)"),
    .INIT(32'h77f344c0))
    al_25e520e0 (
    .a(al_70727c2f),
    .b(al_6aaeddf4),
    .c(al_88fb5330[24]),
    .d(al_a9336f5),
    .e(al_9993ad5e),
    .o(s_axi_rdata[24]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_2fd5aaa (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[25]),
    .d(al_d1b76c6b[25]),
    .e(al_752f7592[25]),
    .o(al_c00b2fb7));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_967da2f6 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[57]),
    .d(al_d1b76c6b[57]),
    .e(al_752f7592[57]),
    .o(al_350ee797));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(~D*B)*~(~E*A))"),
    .INIT(64'h0f030501ff335511))
    al_402e7a72 (
    .a(al_627de329),
    .b(al_fc03cb77),
    .c(al_ce826c89),
    .d(al_c00b2fb7),
    .e(al_350ee797),
    .f(al_49a90ce2[25]),
    .o(al_e5314cad));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))*~(B)+~E*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*~(B)+~(~E)*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*B+~E*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*B)"),
    .INIT(32'h77f344c0))
    al_cef9af15 (
    .a(al_e5314cad),
    .b(al_6aaeddf4),
    .c(al_88fb5330[25]),
    .d(al_a9336f5),
    .e(al_29e11b90),
    .o(s_axi_rdata[25]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_25741d6e (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[26]),
    .d(al_d1b76c6b[26]),
    .e(al_752f7592[26]),
    .o(al_8b041f7e));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_66761479 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[58]),
    .d(al_d1b76c6b[58]),
    .e(al_752f7592[58]),
    .o(al_e5699de4));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(~D*B)*~(~E*A))"),
    .INIT(64'h0f030501ff335511))
    al_92b7ed73 (
    .a(al_627de329),
    .b(al_fc03cb77),
    .c(al_ce826c89),
    .d(al_8b041f7e),
    .e(al_e5699de4),
    .f(al_49a90ce2[26]),
    .o(al_70372a24));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))*~(B)+~E*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*~(B)+~(~E)*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*B+~E*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*B)"),
    .INIT(32'h77f344c0))
    al_508f02a4 (
    .a(al_70372a24),
    .b(al_6aaeddf4),
    .c(al_88fb5330[26]),
    .d(al_a9336f5),
    .e(al_d1a1cb58),
    .o(s_axi_rdata[26]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_3b101d98 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[27]),
    .d(al_d1b76c6b[27]),
    .e(al_752f7592[27]),
    .o(al_87a09a9e));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_31317805 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[59]),
    .d(al_d1b76c6b[59]),
    .e(al_752f7592[59]),
    .o(al_f03a2c10));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(~D*B)*~(~E*A))"),
    .INIT(64'h0f030501ff335511))
    al_80e6ae21 (
    .a(al_627de329),
    .b(al_fc03cb77),
    .c(al_ce826c89),
    .d(al_87a09a9e),
    .e(al_f03a2c10),
    .f(al_49a90ce2[27]),
    .o(al_1824196b));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))*~(B)+~E*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*~(B)+~(~E)*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*B+~E*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*B)"),
    .INIT(32'h77f344c0))
    al_ba7846a6 (
    .a(al_1824196b),
    .b(al_6aaeddf4),
    .c(al_88fb5330[27]),
    .d(al_a9336f5),
    .e(al_989215e7),
    .o(s_axi_rdata[27]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_7c2ea2cc (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[28]),
    .d(al_d1b76c6b[28]),
    .e(al_752f7592[28]),
    .o(al_8765eb4));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_f364a825 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[60]),
    .d(al_d1b76c6b[60]),
    .e(al_752f7592[60]),
    .o(al_3fe33606));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(~D*B)*~(~E*A))"),
    .INIT(64'h0f030501ff335511))
    al_ac9167d (
    .a(al_627de329),
    .b(al_fc03cb77),
    .c(al_ce826c89),
    .d(al_8765eb4),
    .e(al_3fe33606),
    .f(al_49a90ce2[28]),
    .o(al_67074a64));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))*~(B)+~E*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*~(B)+~(~E)*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*B+~E*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*B)"),
    .INIT(32'h77f344c0))
    al_c869b6fc (
    .a(al_67074a64),
    .b(al_6aaeddf4),
    .c(al_88fb5330[28]),
    .d(al_a9336f5),
    .e(al_ac9336a),
    .o(s_axi_rdata[28]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_c52c1fee (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[29]),
    .d(al_d1b76c6b[29]),
    .e(al_752f7592[29]),
    .o(al_9f678f08));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_53bb25a (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[61]),
    .d(al_d1b76c6b[61]),
    .e(al_752f7592[61]),
    .o(al_f6518188));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(~D*B)*~(~E*A))"),
    .INIT(64'h0f030501ff335511))
    al_7c9f1912 (
    .a(al_627de329),
    .b(al_fc03cb77),
    .c(al_ce826c89),
    .d(al_9f678f08),
    .e(al_f6518188),
    .f(al_49a90ce2[29]),
    .o(al_737a8715));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))*~(B)+~E*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*~(B)+~(~E)*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*B+~E*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*B)"),
    .INIT(32'h77f344c0))
    al_b6bb6ae6 (
    .a(al_737a8715),
    .b(al_6aaeddf4),
    .c(al_88fb5330[29]),
    .d(al_a9336f5),
    .e(al_9c616a92),
    .o(s_axi_rdata[29]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_bc1e447d (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[2]),
    .d(al_d1b76c6b[2]),
    .e(al_752f7592[2]),
    .o(al_ff9e33ad));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_81ad05e1 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[34]),
    .d(al_d1b76c6b[34]),
    .e(al_752f7592[34]),
    .o(al_591adfcf));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_5b674f01 (
    .a(al_175588ec),
    .b(al_591adfcf),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_b9297703[2]),
    .f(al_b9297703[3]),
    .o(al_95dcd5c9));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))"),
    .INIT(32'h22200200))
    al_4886a103 (
    .a(al_175588ec),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_49a90ce2[2]),
    .e(al_49a90ce2[34]),
    .o(al_b39aa369));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_3360ded3 (
    .a(al_fc03cb77),
    .b(al_95dcd5c9),
    .c(al_b39aa369),
    .d(al_ff9e33ad),
    .e(al_88fb5330[2]),
    .f(al_a9336f5),
    .o(al_e6b493f[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_4ec127 (
    .a(al_e6b493f[2]),
    .b(al_6aaeddf4),
    .c(al_1974d963),
    .o(s_axi_rdata[2]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*A)"),
    .INIT(64'h0000000000000002))
    al_4fbeb877 (
    .a(s_axi_araddr[7]),
    .b(s_axi_araddr[6]),
    .c(s_axi_araddr[5]),
    .d(s_axi_araddr[4]),
    .e(s_axi_araddr[3]),
    .f(s_axi_araddr[0]),
    .o(al_175588ec));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_1b001734 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[62]),
    .d(al_d1b76c6b[62]),
    .e(al_752f7592[62]),
    .o(al_c2c7d796));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(~D*B)*~(~E*A))"),
    .INIT(64'h0f030501ff335511))
    al_495d2bff (
    .a(al_627de329),
    .b(al_fc03cb77),
    .c(al_ce826c89),
    .d(al_63c928c0),
    .e(al_c2c7d796),
    .f(al_49a90ce2[30]),
    .o(al_90021ccb));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))*~(B)+~E*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*~(B)+~(~E)*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*B+~E*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*B)"),
    .INIT(32'h77f344c0))
    al_144d794 (
    .a(al_90021ccb),
    .b(al_6aaeddf4),
    .c(al_88fb5330[30]),
    .d(al_a9336f5),
    .e(al_e19dcc16),
    .o(s_axi_rdata[30]));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    al_121376ca (
    .a(al_175588ec),
    .b(al_a9336f5),
    .o(al_6aaeddf4));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*B*A)"),
    .INIT(32'h00000080))
    al_1d0192d2 (
    .a(al_175588ec),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_b9297703[2]),
    .e(al_b9297703[3]),
    .o(al_627de329));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~(A*~(~C*B)))"),
    .INIT(32'h0000005d))
    al_a0228cf8 (
    .a(al_175588ec),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_b9297703[2]),
    .e(al_b9297703[3]),
    .o(al_fc03cb77));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_5eb2f895 (
    .a(al_175588ec),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .o(al_ce826c89));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_67414628 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[30]),
    .d(al_d1b76c6b[30]),
    .e(al_752f7592[30]),
    .o(al_63c928c0));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_6308e91b (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[31]),
    .d(al_d1b76c6b[31]),
    .e(al_752f7592[31]),
    .o(al_c58b187c));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_d41b803e (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[63]),
    .d(al_d1b76c6b[63]),
    .e(al_752f7592[63]),
    .o(al_e6bb9c83));
  AL_MAP_LUT6 #(
    .EQN("(~(F*C)*~(~D*B)*~(~E*A))"),
    .INIT(64'h0f030501ff335511))
    al_5905731c (
    .a(al_627de329),
    .b(al_fc03cb77),
    .c(al_ce826c89),
    .d(al_c58b187c),
    .e(al_e6bb9c83),
    .f(al_49a90ce2[31]),
    .o(al_4c4d90b0));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~((~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))*~(B)+~E*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*~(B)+~(~E)*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*B+~E*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)*B)"),
    .INIT(32'h77f344c0))
    al_a7dddc4b (
    .a(al_4c4d90b0),
    .b(al_6aaeddf4),
    .c(al_88fb5330[31]),
    .d(al_a9336f5),
    .e(al_a4c57dd8),
    .o(s_axi_rdata[31]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_d8de005a (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[3]),
    .d(al_d1b76c6b[3]),
    .e(al_752f7592[3]),
    .o(al_a9aea0ae));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_62ed0a48 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[35]),
    .d(al_d1b76c6b[35]),
    .e(al_752f7592[35]),
    .o(al_7a5b596f));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_65abc412 (
    .a(al_175588ec),
    .b(al_7a5b596f),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_b9297703[2]),
    .f(al_b9297703[3]),
    .o(al_e7f17f52));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))"),
    .INIT(32'h22200200))
    al_d9a19ad8 (
    .a(al_175588ec),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_49a90ce2[3]),
    .e(al_49a90ce2[35]),
    .o(al_60993b86));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_d9e939be (
    .a(al_fc03cb77),
    .b(al_e7f17f52),
    .c(al_60993b86),
    .d(al_a9aea0ae),
    .e(al_88fb5330[3]),
    .f(al_a9336f5),
    .o(al_e6b493f[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_ee218db9 (
    .a(al_e6b493f[3]),
    .b(al_6aaeddf4),
    .c(al_b3009928),
    .o(s_axi_rdata[3]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_e90e52e6 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[4]),
    .d(al_d1b76c6b[4]),
    .e(al_752f7592[4]),
    .o(al_ae33357f));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_66391a04 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[36]),
    .d(al_d1b76c6b[36]),
    .e(al_752f7592[36]),
    .o(al_67b92cd9));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_85530a18 (
    .a(al_175588ec),
    .b(al_67b92cd9),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_b9297703[2]),
    .f(al_b9297703[3]),
    .o(al_e774f130));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))"),
    .INIT(32'h22200200))
    al_8fcad573 (
    .a(al_175588ec),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_49a90ce2[4]),
    .e(al_49a90ce2[36]),
    .o(al_edca2c86));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_ad7985cf (
    .a(al_fc03cb77),
    .b(al_e774f130),
    .c(al_edca2c86),
    .d(al_ae33357f),
    .e(al_88fb5330[4]),
    .f(al_a9336f5),
    .o(al_e6b493f[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_1920717d (
    .a(al_e6b493f[4]),
    .b(al_6aaeddf4),
    .c(al_f13bd74f),
    .o(s_axi_rdata[4]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_4b7b4b9d (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[5]),
    .d(al_d1b76c6b[5]),
    .e(al_752f7592[5]),
    .o(al_a7af4189));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_1c64788b (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[37]),
    .d(al_d1b76c6b[37]),
    .e(al_752f7592[37]),
    .o(al_32667361));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_7fd5cea2 (
    .a(al_175588ec),
    .b(al_32667361),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_b9297703[2]),
    .f(al_b9297703[3]),
    .o(al_7ce61a6c));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))"),
    .INIT(32'h22200200))
    al_a7021d8c (
    .a(al_175588ec),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_49a90ce2[5]),
    .e(al_49a90ce2[37]),
    .o(al_711d3f5));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_730dcc (
    .a(al_fc03cb77),
    .b(al_7ce61a6c),
    .c(al_711d3f5),
    .d(al_a7af4189),
    .e(al_88fb5330[5]),
    .f(al_a9336f5),
    .o(al_e6b493f[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_9a188e10 (
    .a(al_e6b493f[5]),
    .b(al_6aaeddf4),
    .c(al_2ad06c7e),
    .o(s_axi_rdata[5]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_d5e607b (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[6]),
    .d(al_d1b76c6b[6]),
    .e(al_752f7592[6]),
    .o(al_2e8c1b28));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_907aa90e (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[38]),
    .d(al_d1b76c6b[38]),
    .e(al_752f7592[38]),
    .o(al_68258153));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_d1a144d3 (
    .a(al_175588ec),
    .b(al_68258153),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_b9297703[2]),
    .f(al_b9297703[3]),
    .o(al_b292fc1));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))"),
    .INIT(32'h22200200))
    al_f8753106 (
    .a(al_175588ec),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_49a90ce2[6]),
    .e(al_49a90ce2[38]),
    .o(al_3c3908e6));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_f807612b (
    .a(al_fc03cb77),
    .b(al_b292fc1),
    .c(al_3c3908e6),
    .d(al_2e8c1b28),
    .e(al_88fb5330[6]),
    .f(al_a9336f5),
    .o(al_e6b493f[6]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_6d6096e (
    .a(al_e6b493f[6]),
    .b(al_6aaeddf4),
    .c(al_159c9d41),
    .o(s_axi_rdata[6]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_6fc56f09 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[7]),
    .d(al_d1b76c6b[7]),
    .e(al_752f7592[7]),
    .o(al_438ac6ff));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_a6804370 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[39]),
    .d(al_d1b76c6b[39]),
    .e(al_752f7592[39]),
    .o(al_ca04b07a));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_adf36d6b (
    .a(al_175588ec),
    .b(al_ca04b07a),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_b9297703[2]),
    .f(al_b9297703[3]),
    .o(al_9e1e2a36));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))"),
    .INIT(32'h22200200))
    al_6b1454d1 (
    .a(al_175588ec),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_49a90ce2[7]),
    .e(al_49a90ce2[39]),
    .o(al_da959817));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_1aa78c58 (
    .a(al_fc03cb77),
    .b(al_9e1e2a36),
    .c(al_da959817),
    .d(al_438ac6ff),
    .e(al_88fb5330[7]),
    .f(al_a9336f5),
    .o(al_e6b493f[7]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_e65f41e (
    .a(al_e6b493f[7]),
    .b(al_6aaeddf4),
    .c(al_fefd5fd3),
    .o(s_axi_rdata[7]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_ef58fb82 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[8]),
    .d(al_d1b76c6b[8]),
    .e(al_752f7592[8]),
    .o(al_da9cd0a9));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_c152d923 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[40]),
    .d(al_d1b76c6b[40]),
    .e(al_752f7592[40]),
    .o(al_d8bac65b));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_f6b1a038 (
    .a(al_175588ec),
    .b(al_d8bac65b),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_b9297703[2]),
    .f(al_b9297703[3]),
    .o(al_8fcbb835));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))"),
    .INIT(32'h22200200))
    al_bf88b32e (
    .a(al_175588ec),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_49a90ce2[8]),
    .e(al_49a90ce2[40]),
    .o(al_ef45b73e));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_e0b7082a (
    .a(al_fc03cb77),
    .b(al_8fcbb835),
    .c(al_ef45b73e),
    .d(al_da9cd0a9),
    .e(al_88fb5330[8]),
    .f(al_a9336f5),
    .o(al_e6b493f[8]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_bf79599a (
    .a(al_e6b493f[8]),
    .b(al_6aaeddf4),
    .c(al_ca969cfa),
    .o(s_axi_rdata[8]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_176d6253 (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[9]),
    .d(al_d1b76c6b[9]),
    .e(al_752f7592[9]),
    .o(al_2c95779d));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8cae9dbf))
    al_ae98b70b (
    .a(al_b9297703[0]),
    .b(al_b9297703[1]),
    .c(al_902efd00[41]),
    .d(al_d1b76c6b[41]),
    .e(al_752f7592[41]),
    .o(al_edb0b8cc));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*~B*A)"),
    .INIT(64'h0000000000002000))
    al_f51b1254 (
    .a(al_175588ec),
    .b(al_edb0b8cc),
    .c(s_axi_araddr[2]),
    .d(s_axi_araddr[1]),
    .e(al_b9297703[2]),
    .f(al_b9297703[3]),
    .o(al_6e6c13e6));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))"),
    .INIT(32'h22200200))
    al_cdd3b8f2 (
    .a(al_175588ec),
    .b(s_axi_araddr[2]),
    .c(s_axi_araddr[1]),
    .d(al_49a90ce2[9]),
    .e(al_49a90ce2[41]),
    .o(al_f7e49aaa));
  AL_MAP_LUT6 #(
    .EQN("~(~E*~((~C*~B*~(~D*A)))*~(F)+~E*(~C*~B*~(~D*A))*~(F)+~(~E)*(~C*~B*~(~D*A))*F+~E*(~C*~B*~(~D*A))*F)"),
    .INIT(64'hfcfefcfeffff0000))
    al_526d020c (
    .a(al_fc03cb77),
    .b(al_6e6c13e6),
    .c(al_f7e49aaa),
    .d(al_2c95779d),
    .e(al_88fb5330[9]),
    .f(al_a9336f5),
    .o(al_e6b493f[9]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_563204a8 (
    .a(al_e6b493f[9]),
    .b(al_6aaeddf4),
    .c(al_dd993167),
    .o(s_axi_rdata[9]));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    al_9e8e6d55 (
    .a(al_6ea32e9c),
    .o(speed_1000));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_817c9c10 (
    .a(speed_100),
    .b(al_6ea32e9c),
    .o(speed_10));

endmodule 

